
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_FPmul is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_FPmul;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         FP_Z : out std_logic_vector (31 downto 0));

end FPmul;

architecture SYN_pipeline of FPmul is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal A_EXP_7_port, A_EXP_6_port, A_EXP_5_port, A_EXP_4_port, A_EXP_3_port,
      A_EXP_2_port, A_EXP_1_port, A_EXP_0_port, A_SIG_8_port, B_EXP_7_port, 
      B_EXP_6_port, B_EXP_5_port, B_EXP_4_port, B_EXP_3_port, B_EXP_2_port, 
      B_EXP_1_port, B_EXP_0_port, B_SIG_9_port, B_SIG_8_port, SIGN_out_stage1, 
      isINF_stage1, isNaN_stage1, isZ_tab_stage1, EXP_in_7_port, EXP_in_3_port,
      EXP_in_2_port, EXP_neg_stage2, EXP_pos_stage2, SIGN_out_stage2, 
      SIG_in_27_port, isINF_stage2, isNaN_stage2, isZ_tab_stage2, EXP_neg, 
      EXP_out_round_7_port, EXP_out_round_4_port, EXP_out_round_3_port, 
      EXP_out_round_2_port, EXP_out_round_1_port, I1_isZ_tab_int, I1_isNaN_int,
      I1_isINF_int, I1_SIGN_out_int, I2_dtemp_30_port, I2_dtemp_31_port, 
      I2_dtemp_33_port, I2_dtemp_34_port, I2_dtemp_39_port, I2_dtemp_41_port, 
      I2_dtemp_42_port, I2_dtemp_43_port, I2_dtemp_44_port, I2_mw_I4sum_0_port,
      I2_mw_I4sum_1_port, I2_mw_I4sum_2_port, I2_mw_I4sum_3_port, 
      I2_mw_I4sum_4_port, I2_mw_I4sum_5_port, I2_mw_I4sum_6_port, I2_N0, 
      I2_SIGN_out_stage2_tmp, I2_isZ_tab_stage2_tmp, I2_isNaN_stage2_tmp, 
      I2_isINF_stage2_tmp, I2_EXP_neg_stage2_tmp, I2_EXP_pos_int, 
      I2_EXP_pos_stage2_tmp, I2_EXP_in_tmp_0_port, I2_EXP_in_tmp_1_port, 
      I2_EXP_in_tmp_2_port, I2_EXP_in_tmp_3_port, I2_EXP_in_tmp_5_port, 
      I2_EXP_in_tmp_6_port, I2_EXP_in_tmp_7_port, I3_SIG_out_4_port, 
      I3_SIG_out_5_port, I3_SIG_out_6_port, I3_SIG_out_7_port, 
      I3_SIG_out_8_port, I3_SIG_out_9_port, I3_SIG_out_10_port, 
      I3_SIG_out_11_port, I3_SIG_out_12_port, I3_SIG_out_13_port, 
      I3_SIG_out_14_port, I3_SIG_out_15_port, I3_SIG_out_16_port, 
      I3_SIG_out_17_port, I3_SIG_out_18_port, I3_SIG_out_19_port, 
      I3_EXP_out_0_port, I3_EXP_out_1_port, I3_EXP_out_2_port, 
      I3_EXP_out_3_port, I3_EXP_out_4_port, I3_EXP_out_5_port, 
      I3_EXP_out_6_port, I3_EXP_out_7_port, I4_FP_31_port, I1_I0_N13, I1_I1_N13
      , n359, n360, n374, n381, n384, n2556, n2557, n2558, n2559, n2560, n2561,
      n2562, n2563, n2565, n2567, n2568, n2569, n2570, n2571, n2572, n2573, 
      n2574, n2577, n2579, n2583, n2584, n2587, n2589, n2590, n2592, n2593, 
      n2594, n2596, n2597, n2598, n2602, n2606, n2611, n2613, n2638, n4381, 
      n8323, n8325, n8326, n8329, n8330, n8331, n8332, n8333, n8334, n8338, 
      n8339, n8340, n8345, n8346, n8347, n8349, n8350, n8351, n8352, n8353, 
      n8355, n8358, n8363, n8371, n8374, n8375, n8376, n8379, n8381, n8385, 
      n8391, n8392, n8401, n8406, n8409, n10593, n10596, intadd_42_A_3_port, 
      intadd_42_B_3_port, intadd_42_n11, intadd_56_A_3_port, intadd_66_A_1_port
      , intadd_66_A_0_port, intadd_66_B_1_port, intadd_66_B_0_port, 
      intadd_66_CI, intadd_66_SUM_2_port, intadd_66_SUM_1_port, intadd_66_n3, 
      intadd_66_n2, intadd_66_n1, intadd_47_SUM_3_port, intadd_46_A_3_port, 
      intadd_46_A_2_port, intadd_46_A_1_port, intadd_46_B_4_port, 
      intadd_46_B_3_port, intadd_46_B_1_port, intadd_46_B_0_port, intadd_46_CI,
      intadd_46_SUM_4_port, intadd_46_SUM_3_port, intadd_46_SUM_2_port, 
      intadd_46_SUM_1_port, intadd_46_SUM_0_port, intadd_46_n5, intadd_46_n4, 
      intadd_46_n3, intadd_46_n2, intadd_46_n1, intadd_58_A_2_port, 
      intadd_58_A_1_port, intadd_58_A_0_port, intadd_58_B_2_port, 
      intadd_58_B_1_port, intadd_58_B_0_port, intadd_58_CI, 
      intadd_58_SUM_2_port, intadd_58_SUM_1_port, intadd_58_SUM_0_port, 
      intadd_58_n3, intadd_58_n2, intadd_58_n1, intadd_62_A_2_port, 
      intadd_62_A_1_port, intadd_62_A_0_port, intadd_62_B_2_port, 
      intadd_62_B_1_port, intadd_62_B_0_port, intadd_62_CI, 
      intadd_62_SUM_2_port, intadd_62_SUM_1_port, intadd_62_SUM_0_port, 
      intadd_62_n3, intadd_62_n2, intadd_62_n1, intadd_61_n7, intadd_61_n6, 
      intadd_61_n5, intadd_61_n2, intadd_61_n1, intadd_63_SUM_2_port, n10597, 
      n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10607, 
      n10608, n10609, n10610, n10611, n10613, n10614, n10615, n10617, n10618, 
      n10619, n10620, n10621, n10623, n10624, n10625, n10626, n10627, n10630, 
      n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, 
      n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, 
      n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, 
      n10658, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, 
      n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, 
      n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, 
      n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, 
      n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, 
      n10705, n10707, n10708, n10709, n10710, n10711, n10713, n10714, n10715, 
      n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, 
      n10725, n10726, n10727, n10728, n10730, n10731, n10733, n10734, n10736, 
      n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, 
      n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, 
      n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, 
      n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, 
      n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, 
      n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, 
      n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, 
      n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, 
      n10809, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, 
      n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, 
      n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, 
      n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, 
      n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, 
      n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, 
      n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, 
      n10873, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, 
      n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, 
      n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, 
      n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, 
      n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, 
      n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, 
      n10928, n10929, n10930, n10931, n10932, n10934, n10935, n10936, n10937, 
      n10938, n10939, n10940, n10942, n10943, n10944, n10945, n10947, n10948, 
      n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10958, 
      n10959, n10960, n10963, n10964, n10965, n10966, n10967, n10968, n10969, 
      n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, 
      n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, 
      n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, 
      n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, 
      n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, 
      n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, 
      n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, 
      n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, 
      n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, 
      n11051, n11052, n11053, n11054, n11056, n11057, n11058, n11059, n11060, 
      n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, 
      n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, 
      n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, 
      n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, 
      n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, 
      n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, 
      n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, 
      n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, 
      n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, 
      n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, 
      n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, 
      n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, 
      n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, 
      n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, 
      n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, 
      n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, 
      n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, 
      n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, 
      n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, 
      n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, 
      n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, 
      n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, 
      n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, 
      n11269, n11270, n11271, n11272, n11274, n11275, n11276, n11277, n11278, 
      n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, 
      n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, 
      n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, 
      n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, 
      n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11324, 
      n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, 
      n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, 
      n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, 
      n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, 
      n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, 
      n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, 
      n11379, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11389, 
      n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, 
      n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, 
      n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, 
      n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, 
      n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, 
      n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, 
      n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, 
      n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, 
      n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, 
      n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, 
      n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, 
      n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, 
      n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, 
      n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, 
      n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, 
      n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, 
      n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, 
      n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, 
      n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, 
      n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, 
      n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, 
      n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, 
      n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11596, n11597, 
      n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, 
      n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, 
      n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, 
      n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, 
      n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, 
      n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, 
      n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, 
      n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, 
      n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, 
      n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, 
      n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, 
      n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, 
      n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, 
      n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, 
      n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, 
      n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, 
      n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, 
      n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, 
      n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, 
      n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, 
      n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, 
      n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, 
      n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, 
      n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, 
      n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, 
      n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, 
      n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, 
      n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, 
      n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, 
      n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, 
      n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, 
      n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, 
      n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, 
      n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, 
      n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, 
      n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, 
      n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, 
      n11931, n11932, n11933, n11935, n11936, n11937, n11938, n11939, n11940, 
      n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, 
      n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, 
      n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, 
      n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, 
      n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, 
      n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, 
      n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, 
      n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, 
      n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, 
      n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, 
      n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12040, 
      n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, 
      n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, 
      n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, 
      n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, 
      n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, 
      n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, 
      n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, 
      n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, 
      n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, 
      n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, 
      n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, 
      n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, 
      n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, 
      n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, 
      n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, 
      n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, 
      n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, 
      n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, 
      n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, 
      n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, 
      n12221, n12222, n12223, n12224, n12225, n12226, n12228, n12229, n12230, 
      n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, 
      n12240, n12241, n12243, n12244, n12245, n12246, n12247, n12248, n12249, 
      n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, 
      n12259, n12260, n12261, n12262, n12264, n12265, n12267, n12268, n12269, 
      n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, 
      n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, 
      n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, 
      n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, 
      n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, 
      n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, 
      n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, 
      n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, 
      n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, 
      n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, 
      n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, 
      n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, 
      n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, 
      n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, 
      n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, 
      n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, 
      n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, 
      n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, 
      n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, 
      n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, 
      n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, 
      n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, 
      n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, 
      n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, 
      n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, 
      n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, 
      n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, 
      n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, 
      n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, 
      n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, 
      n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, 
      n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, 
      n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, 
      n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, 
      n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, 
      n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, 
      n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, 
      n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, 
      n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, 
      n12623, n12624, n12625, n12627, n12628, n12629, n12630, n12631, n12632, 
      n12633, n12634, n12636, n12637, n12638, n12639, n12640, n12641, n12642, 
      n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, 
      n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, 
      n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, 
      n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, 
      n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, 
      n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, 
      n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, 
      n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, 
      n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, 
      n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, 
      n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, 
      n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, 
      n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, 
      n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, 
      n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, 
      n12778, n12779, n12780, n12781, n12782, n12783, n12785, n12786, n12787, 
      n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, 
      n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, 
      n12806, n12807, n12808, n12809, n12811, n12812, n12813, n12814, n12815, 
      n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, 
      n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, 
      n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, 
      n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, 
      n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, 
      n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, 
      n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, 
      n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, 
      n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, 
      n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, 
      n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, 
      n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, 
      n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, 
      n12933, n12934, n12935, n12937, n12938, n12939, n12940, n12941, n12942, 
      n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, 
      n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, 
      n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, 
      n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, 
      n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, 
      n12988, n12989, n12990, n12992, n12993, n12994, n12995, n12996, n12997, 
      n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, 
      n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, 
      n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, 
      n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, 
      n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, 
      n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, 
      n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, 
      n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, 
      n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, 
      n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, 
      n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, 
      n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, 
      n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, 
      n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, 
      n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, 
      n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, 
      n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, 
      n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, 
      n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, 
      n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13177, n13178, 
      n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, 
      n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, 
      n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, 
      n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, 
      n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, 
      n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, 
      n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, 
      n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, 
      n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, 
      n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, 
      n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, 
      n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, 
      n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, 
      n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, 
      n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, 
      n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, 
      n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, 
      n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, 
      n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, 
      n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, 
      n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, 
      n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, 
      n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, 
      n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, 
      n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, 
      n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, 
      n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, 
      n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, 
      n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, 
      n13440, n13442, n13443, n13444, n13445, n13447, n13448, n13449, n13450, 
      n13451, n13452, n13453, n13454, n13456, n13457, n13458, n13459, n13460, 
      n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, 
      n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, 
      n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, 
      n13488, n13489, n13490, n13491, n13492, n13493, n13495, n13496, n13497, 
      n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, 
      n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, 
      n13516, n13517, n13518, n13520, n13521, n13522, n13523, n13524, n13525, 
      n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, 
      n13535, n13536, n13537, n13538, n13539, n13540, n13542, n13543, n13544, 
      n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, 
      n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, 
      n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, 
      n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, 
      n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, 
      n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, 
      n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, 
      n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, 
      n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, 
      n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, 
      n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, 
      n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, 
      n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, 
      n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, 
      n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, 
      n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, 
      n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, 
      n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, 
      n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, 
      n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, 
      n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, 
      n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, 
      n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, 
      n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, 
      n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, 
      n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, 
      n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, 
      n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, 
      n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, 
      n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, 
      n13816, n13817, n13819, n13820, n13821, n13822, n13823, n13824, n13825, 
      n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, 
      n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, 
      n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, 
      n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, 
      n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, 
      n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, 
      n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, 
      n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, 
      n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, 
      n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, 
      n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, 
      n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, 
      n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, 
      n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, 
      n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, 
      n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, 
      n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, 
      n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, 
      n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, 
      n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, 
      n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, 
      n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, 
      n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, 
      n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, 
      n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, 
      n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, 
      n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, 
      n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, 
      n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, 
      n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, 
      n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, 
      n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, 
      n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, 
      n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, 
      n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, 
      n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, 
      n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, 
      n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, 
      n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, 
      n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, 
      n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, 
      n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14205, 
      n14206, n14207, n14209, n14210, n14211, n14212, n14213, n14214, n14215, 
      n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, 
      n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, 
      n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, 
      n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, 
      n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, 
      n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, 
      n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, 
      n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, 
      n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, 
      n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, 
      n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, 
      n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, 
      n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, 
      n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, 
      n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, 
      n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, 
      n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, 
      n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, 
      n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, 
      n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, 
      n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, 
      n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, 
      n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, 
      n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, 
      n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, 
      n14441, n14442, n14446, n14447, n14448, n14449, n14450, n14451, n14452, 
      n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, 
      n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, 
      n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, 
      n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, 
      n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, 
      n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, 
      n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, 
      n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, 
      n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, 
      n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, 
      n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, 
      n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, 
      n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, 
      n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, 
      n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, 
      n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, 
      n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, 
      n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, 
      n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, 
      n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, 
      n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, 
      n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, 
      n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, 
      n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, 
      n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, 
      n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, 
      n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, 
      n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, 
      n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, 
      n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, 
      n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, 
      n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, 
      n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, 
      n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, 
      n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, 
      n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, 
      n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, 
      n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, 
      n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, 
      n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, 
      n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, 
      n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, 
      n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, 
      n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, 
      n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, 
      n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, 
      n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, 
      n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, 
      n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, 
      n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, 
      n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, 
      n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, 
      n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, 
      n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14940, 
      n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, 
      n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, 
      n14959, n14960, n14961, n14962, n14963, n14964, n14965, n_1000, n_1001, 
      n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, 
      n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, 
      n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, 
      n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, 
      n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, 
      n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, 
      n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, 
      n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, 
      n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, 
      n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, 
      n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, 
      n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, 
      n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, 
      n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, 
      n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, 
      n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, 
      n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, 
      n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, 
      n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, 
      n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, 
      n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, 
      n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, 
      n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, 
      n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, 
      n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, 
      n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, 
      n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, 
      n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, 
      n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, 
      n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, 
      n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, 
      n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, 
      n_1353, n_1354 : std_logic;

begin
   
   I1_B_EXP_reg_0_inst : DFF_X1 port map( D => FP_B(23), CK => clk, Q => 
                           B_EXP_0_port, QN => n_1000);
   I1_B_EXP_reg_1_inst : DFF_X1 port map( D => FP_B(24), CK => clk, Q => 
                           B_EXP_1_port, QN => n_1001);
   I1_B_EXP_reg_4_inst : DFF_X1 port map( D => FP_B(27), CK => clk, Q => 
                           B_EXP_4_port, QN => n14475);
   I1_B_EXP_reg_5_inst : DFF_X1 port map( D => FP_B(28), CK => clk, Q => 
                           B_EXP_5_port, QN => n_1002);
   I1_B_EXP_reg_6_inst : DFF_X1 port map( D => FP_B(29), CK => clk, Q => 
                           B_EXP_6_port, QN => n14474);
   I1_B_EXP_reg_7_inst : DFF_X1 port map( D => FP_B(30), CK => clk, Q => 
                           B_EXP_7_port, QN => n_1003);
   I1_isNaN_stage1_reg : DFF_X1 port map( D => I1_isNaN_int, CK => clk, Q => 
                           isNaN_stage1, QN => n_1004);
   I1_isINF_stage1_reg : DFF_X1 port map( D => I1_isINF_int, CK => clk, Q => 
                           isINF_stage1, QN => n_1005);
   R_1460 : DFF_X1 port map( D => FP_A(4), CK => clk, Q => n8363, QN => n10639)
                           ;
   R_1286 : DFF_X1 port map( D => FP_A(6), CK => clk, Q => n_1006, QN => n14597
                           );
   R_1515 : DFF_X1 port map( D => FP_A(10), CK => clk, Q => n14488, QN => 
                           n_1007);
   R_1327 : DFF_X1 port map( D => FP_A(12), CK => clk, Q => n10690, QN => 
                           n14584);
   R_1457 : DFF_X1 port map( D => FP_A(14), CK => clk, Q => n_1008, QN => 
                           n10884);
   R_0 : DFF_X1 port map( D => FP_A(18), CK => clk, Q => n10935, QN => n14711);
   I1_A_EXP_reg_0_inst : DFF_X1 port map( D => FP_A(23), CK => clk, Q => 
                           A_EXP_0_port, QN => n_1009);
   I1_A_EXP_reg_1_inst : DFF_X1 port map( D => FP_A(24), CK => clk, Q => 
                           A_EXP_1_port, QN => n_1010);
   I1_A_EXP_reg_3_inst : DFF_X1 port map( D => FP_A(26), CK => clk, Q => 
                           A_EXP_3_port, QN => n14504);
   I1_A_EXP_reg_4_inst : DFF_X1 port map( D => FP_A(27), CK => clk, Q => 
                           A_EXP_4_port, QN => n14506);
   I1_A_EXP_reg_5_inst : DFF_X1 port map( D => FP_A(28), CK => clk, Q => 
                           A_EXP_5_port, QN => n_1011);
   I1_A_EXP_reg_6_inst : DFF_X1 port map( D => FP_A(29), CK => clk, Q => 
                           A_EXP_6_port, QN => n14503);
   I1_A_EXP_reg_7_inst : DFF_X1 port map( D => FP_A(30), CK => clk, Q => 
                           A_EXP_7_port, QN => n_1012);
   I1_SIGN_out_stage1_reg : DFF_X1 port map( D => I1_SIGN_out_int, CK => clk, Q
                           => SIGN_out_stage1, QN => n_1013);
   I2_SIGN_out_stage2_tmp_reg : DFF_X1 port map( D => SIGN_out_stage1, CK => 
                           clk, Q => I2_SIGN_out_stage2_tmp, QN => n_1014);
   I2_SIGN_out_stage2_reg : DFF_X1 port map( D => I2_SIGN_out_stage2_tmp, CK =>
                           clk, Q => SIGN_out_stage2, QN => n_1015);
   I2_isZ_tab_stage2_tmp_reg : DFF_X1 port map( D => isZ_tab_stage1, CK => clk,
                           Q => I2_isZ_tab_stage2_tmp, QN => n_1016);
   I2_isZ_tab_stage2_reg : DFF_X1 port map( D => I2_isZ_tab_stage2_tmp, CK => 
                           clk, Q => isZ_tab_stage2, QN => n_1017);
   I2_isNaN_stage2_tmp_reg : DFF_X1 port map( D => isNaN_stage1, CK => clk, Q 
                           => I2_isNaN_stage2_tmp, QN => n_1018);
   I2_isNaN_stage2_reg : DFF_X1 port map( D => I2_isNaN_stage2_tmp, CK => clk, 
                           Q => isNaN_stage2, QN => n_1019);
   I2_isINF_stage2_tmp_reg : DFF_X1 port map( D => isINF_stage1, CK => clk, Q 
                           => I2_isINF_stage2_tmp, QN => n_1020);
   I2_isINF_stage2_reg : DFF_X1 port map( D => I2_isINF_stage2_tmp, CK => clk, 
                           Q => isINF_stage2, QN => n_1021);
   I2_EXP_neg_stage2_tmp_reg : DFF_X1 port map( D => I2_N0, CK => clk, Q => 
                           I2_EXP_neg_stage2_tmp, QN => n_1022);
   I2_EXP_neg_stage2_reg : DFF_X1 port map( D => I2_EXP_neg_stage2_tmp, CK => 
                           clk, Q => EXP_neg_stage2, QN => n_1023);
   I2_EXP_pos_stage2_tmp_reg : DFF_X1 port map( D => I2_EXP_pos_int, CK => clk,
                           Q => I2_EXP_pos_stage2_tmp, QN => n_1024);
   I2_EXP_pos_stage2_reg : DFF_X1 port map( D => I2_EXP_pos_stage2_tmp, CK => 
                           clk, Q => EXP_pos_stage2, QN => n_1025);
   R_1333 : DFF_X1 port map( D => n14490, CK => clk, Q => n10943, QN => n_1026)
                           ;
   I2_SIG_in_reg_8_inst : DFF_X1 port map( D => n14517, CK => clk, Q => n14471,
                           QN => n2606);
   I2_SIG_in_reg_9_inst : DFF_X1 port map( D => n8406, CK => clk, Q => n8381, 
                           QN => n14519);
   I2_SIG_in_reg_10_inst : DFF_X1 port map( D => I2_dtemp_30_port, CK => clk, Q
                           => n8371, QN => n_1027);
   I2_SIG_in_reg_12_inst : DFF_X1 port map( D => n10593, CK => clk, Q => n_1028
                           , QN => n2602);
   I2_SIG_in_reg_14_inst : DFF_X1 port map( D => I2_dtemp_34_port, CK => clk, Q
                           => n14497, QN => n_1029);
   I2_SIG_in_reg_15_inst : DFF_X1 port map( D => n14937, CK => clk, Q => n8346,
                           QN => n_1030);
   I2_SIG_in_reg_17_inst : DFF_X1 port map( D => n14933, CK => clk, Q => n_1031
                           , QN => n2597);
   I2_SIG_in_reg_24_inst : DFF_X1 port map( D => I2_dtemp_44_port, CK => clk, Q
                           => n_1032, QN => n2590);
   I2_EXP_in_tmp_reg_0_inst : DFF_X1 port map( D => I2_mw_I4sum_0_port, CK => 
                           clk, Q => I2_EXP_in_tmp_0_port, QN => n_1033);
   I2_EXP_in_tmp_reg_1_inst : DFF_X1 port map( D => I2_mw_I4sum_1_port, CK => 
                           clk, Q => I2_EXP_in_tmp_1_port, QN => n_1034);
   I2_EXP_in_reg_1_inst : DFF_X1 port map( D => I2_EXP_in_tmp_1_port, CK => clk
                           , Q => n_1035, QN => n2577);
   I2_EXP_in_tmp_reg_2_inst : DFF_X1 port map( D => I2_mw_I4sum_2_port, CK => 
                           clk, Q => I2_EXP_in_tmp_2_port, QN => n_1036);
   I2_EXP_in_tmp_reg_3_inst : DFF_X1 port map( D => I2_mw_I4sum_3_port, CK => 
                           clk, Q => I2_EXP_in_tmp_3_port, QN => n_1037);
   I2_EXP_in_reg_3_inst : DFF_X1 port map( D => I2_EXP_in_tmp_3_port, CK => clk
                           , Q => EXP_in_3_port, QN => n14511);
   I2_EXP_in_tmp_reg_5_inst : DFF_X1 port map( D => I2_mw_I4sum_5_port, CK => 
                           clk, Q => I2_EXP_in_tmp_5_port, QN => n_1038);
   I2_EXP_in_reg_5_inst : DFF_X1 port map( D => I2_EXP_in_tmp_5_port, CK => clk
                           , Q => n_1039, QN => n14493);
   I2_EXP_in_tmp_reg_6_inst : DFF_X1 port map( D => I2_mw_I4sum_6_port, CK => 
                           clk, Q => I2_EXP_in_tmp_6_port, QN => n_1040);
   I2_EXP_in_tmp_reg_7_inst : DFF_X1 port map( D => n374, CK => clk, Q => 
                           I2_EXP_in_tmp_7_port, QN => n_1041);
   I2_EXP_in_reg_7_inst : DFF_X1 port map( D => I2_EXP_in_tmp_7_port, CK => clk
                           , Q => EXP_in_7_port, QN => n_1042);
   I3_EXP_neg_reg : DFF_X1 port map( D => EXP_neg_stage2, CK => clk, Q => 
                           EXP_neg, QN => n_1043);
   I3_EXP_pos_reg : DFF_X1 port map( D => EXP_pos_stage2, CK => clk, Q => 
                           n_1044, QN => n2613);
   I3_SIGN_out_reg : DFF_X1 port map( D => SIGN_out_stage2, CK => clk, Q => 
                           I4_FP_31_port, QN => n_1045);
   I3_isZ_tab_reg : DFF_X1 port map( D => isZ_tab_stage2, CK => clk, Q => 
                           n_1046, QN => n2611);
   I3_isNaN_reg : DFF_X1 port map( D => isNaN_stage2, CK => clk, Q => n_1047, 
                           QN => n2567);
   I3_isINF_tab_reg : DFF_X1 port map( D => isINF_stage2, CK => clk, Q => 
                           n_1048, QN => n8385);
   I3_SIG_out_round_reg_3_inst : DFF_X1 port map( D => n10596, CK => clk, Q => 
                           n_1049, QN => n2587);
   I3_SIG_out_round_reg_4_inst : DFF_X1 port map( D => I3_SIG_out_4_port, CK =>
                           clk, Q => n_1050, QN => n2565);
   I3_SIG_out_round_reg_5_inst : DFF_X1 port map( D => I3_SIG_out_5_port, CK =>
                           clk, Q => n_1051, QN => n2556);
   I3_SIG_out_round_reg_6_inst : DFF_X1 port map( D => I3_SIG_out_6_port, CK =>
                           clk, Q => n_1052, QN => n2568);
   I3_SIG_out_round_reg_7_inst : DFF_X1 port map( D => I3_SIG_out_7_port, CK =>
                           clk, Q => n_1053, QN => n2557);
   I3_SIG_out_round_reg_8_inst : DFF_X1 port map( D => I3_SIG_out_8_port, CK =>
                           clk, Q => n_1054, QN => n2569);
   I3_SIG_out_round_reg_9_inst : DFF_X1 port map( D => I3_SIG_out_9_port, CK =>
                           clk, Q => n_1055, QN => n2558);
   I3_SIG_out_round_reg_10_inst : DFF_X1 port map( D => I3_SIG_out_10_port, CK 
                           => clk, Q => n_1056, QN => n2570);
   I3_SIG_out_round_reg_11_inst : DFF_X1 port map( D => I3_SIG_out_11_port, CK 
                           => clk, Q => n_1057, QN => n2559);
   I3_SIG_out_round_reg_12_inst : DFF_X1 port map( D => I3_SIG_out_12_port, CK 
                           => clk, Q => n_1058, QN => n2571);
   I3_SIG_out_round_reg_13_inst : DFF_X1 port map( D => I3_SIG_out_13_port, CK 
                           => clk, Q => n_1059, QN => n2560);
   I3_SIG_out_round_reg_14_inst : DFF_X1 port map( D => I3_SIG_out_14_port, CK 
                           => clk, Q => n_1060, QN => n2572);
   I3_SIG_out_round_reg_15_inst : DFF_X1 port map( D => I3_SIG_out_15_port, CK 
                           => clk, Q => n_1061, QN => n2561);
   I3_SIG_out_round_reg_16_inst : DFF_X1 port map( D => I3_SIG_out_16_port, CK 
                           => clk, Q => n_1062, QN => n2573);
   I3_SIG_out_round_reg_17_inst : DFF_X1 port map( D => I3_SIG_out_17_port, CK 
                           => clk, Q => n_1063, QN => n2562);
   I3_SIG_out_round_reg_18_inst : DFF_X1 port map( D => I3_SIG_out_18_port, CK 
                           => clk, Q => n_1064, QN => n2574);
   I3_SIG_out_round_reg_19_inst : DFF_X1 port map( D => I3_SIG_out_19_port, CK 
                           => clk, Q => n_1065, QN => n2563);
   I3_EXP_out_round_reg_0_inst : DFF_X1 port map( D => I3_EXP_out_0_port, CK =>
                           clk, Q => n_1066, QN => n2584);
   I3_EXP_out_round_reg_1_inst : DFF_X1 port map( D => I3_EXP_out_1_port, CK =>
                           clk, Q => EXP_out_round_1_port, QN => n_1067);
   I3_EXP_out_round_reg_2_inst : DFF_X1 port map( D => I3_EXP_out_2_port, CK =>
                           clk, Q => EXP_out_round_2_port, QN => n14476);
   I3_EXP_out_round_reg_3_inst : DFF_X1 port map( D => I3_EXP_out_3_port, CK =>
                           clk, Q => EXP_out_round_3_port, QN => n14508);
   I3_EXP_out_round_reg_6_inst : DFF_X1 port map( D => I3_EXP_out_6_port, CK =>
                           clk, Q => n_1068, QN => n2579);
   I4_FP_Z_reg_31_inst : DFF_X1 port map( D => I4_FP_31_port, CK => clk, Q => 
                           FP_Z(31), QN => n_1069);
   I1_isZ_tab_stage1_reg : DFF_X1 port map( D => I1_isZ_tab_int, CK => clk, Q 
                           => isZ_tab_stage1, QN => n_1070);
   R_1477 : DFF_X1 port map( D => FP_A(0), CK => clk, Q => n8358, QN => n14501)
                           ;
   I3_EXP_out_round_reg_7_inst : DFF_X1 port map( D => I3_EXP_out_7_port, CK =>
                           clk, Q => EXP_out_round_7_port, QN => n_1071);
   R_1523 : DFF_X1 port map( D => FP_B(11), CK => clk, Q => n8392, QN => n14457
                           );
   I1_B_SIG_reg_17_inst : DFF_X1 port map( D => FP_B(17), CK => clk, Q => n8330
                           , QN => n14482);
   R_1541 : DFF_X1 port map( D => FP_B(9), CK => clk, Q => B_SIG_9_port, QN => 
                           n14453);
   I1_B_SIG_reg_10_inst : DFF_X1 port map( D => FP_B(10), CK => clk, Q => n8351
                           , QN => n14464);
   I2_EXP_in_reg_0_inst : DFF_X1 port map( D => I2_EXP_in_tmp_0_port, CK => clk
                           , Q => n14502, QN => n2583);
   I2_SIG_in_reg_21_inst : DFF_X1 port map( D => I2_dtemp_41_port, CK => clk, Q
                           => n_1072, QN => n2593);
   I2_SIG_in_reg_19_inst : DFF_X1 port map( D => I2_dtemp_39_port, CK => clk, Q
                           => n8391, QN => n_1073);
   I1_B_SIG_reg_21_inst : DFF_X1 port map( D => FP_B(21), CK => clk, Q => n8334
                           , QN => n14467);
   R_1537 : DFF_X1 port map( D => FP_B(19), CK => clk, Q => n8325, QN => n14466
                           );
   R_1567 : DFF_X2 port map( D => FP_B(16), CK => clk, Q => n14478, QN => 
                           n10831);
   I1_B_EXP_reg_3_inst : DFF_X1 port map( D => FP_B(26), CK => clk, Q => 
                           B_EXP_3_port, QN => n14472);
   I2_EXP_in_reg_4_inst : DFF_X1 port map( D => n8323, CK => clk, Q => n_1074, 
                           QN => n14494);
   I1_B_SIG_reg_20_inst : DFF_X1 port map( D => FP_B(20), CK => clk, Q => n8349
                           , QN => n14458);
   R_1453 : DFF_X1 port map( D => FP_B(18), CK => clk, Q => n8329, QN => n14450
                           );
   R_1539 : DFF_X1 port map( D => FP_B(7), CK => clk, Q => n8333, QN => n14451)
                           ;
   I1_B_SIG_reg_15_inst : DFF_X1 port map( D => FP_B(15), CK => clk, Q => n8332
                           , QN => n14452);
   intadd_66_U4 : FA_X1 port map( A => intadd_66_A_0_port, B => 
                           intadd_66_B_0_port, CI => intadd_66_CI, CO => 
                           intadd_66_n3, S => intadd_56_A_3_port);
   intadd_66_U3 : FA_X1 port map( A => intadd_66_A_1_port, B => 
                           intadd_66_B_1_port, CI => intadd_66_n3, CO => 
                           intadd_66_n2, S => intadd_66_SUM_1_port);
   intadd_46_U6 : FA_X1 port map( A => n14489, B => intadd_46_B_0_port, CI => 
                           intadd_46_CI, CO => intadd_46_n5, S => 
                           intadd_46_SUM_0_port);
   intadd_46_U5 : FA_X1 port map( A => intadd_46_B_1_port, B => 
                           intadd_46_A_1_port, CI => intadd_46_n5, CO => 
                           intadd_46_n4, S => intadd_46_SUM_1_port);
   intadd_46_U4 : FA_X1 port map( A => intadd_46_A_2_port, B => intadd_46_n4, 
                           CI => n14936, CO => intadd_46_n3, S => 
                           intadd_46_SUM_2_port);
   intadd_58_U4 : FA_X1 port map( A => intadd_58_A_0_port, B => 
                           intadd_58_B_0_port, CI => intadd_58_CI, CO => 
                           intadd_58_n3, S => intadd_58_SUM_0_port);
   intadd_58_U3 : FA_X1 port map( A => intadd_58_A_1_port, B => 
                           intadd_58_B_1_port, CI => intadd_58_n3, CO => 
                           intadd_58_n2, S => intadd_58_SUM_1_port);
   intadd_58_U2 : FA_X1 port map( A => intadd_58_A_2_port, B => intadd_58_n2, 
                           CI => intadd_58_B_2_port, CO => intadd_58_n1, S => 
                           intadd_58_SUM_2_port);
   R_1553 : DFF_X1 port map( D => FP_B(4), CK => clk, Q => n8350, QN => n14465)
                           ;
   intadd_62_U4 : FA_X1 port map( A => intadd_62_A_0_port, B => 
                           intadd_62_B_0_port, CI => intadd_62_CI, CO => 
                           intadd_62_n3, S => intadd_62_SUM_0_port);
   intadd_62_U3 : FA_X1 port map( A => intadd_62_A_1_port, B => 
                           intadd_62_B_1_port, CI => intadd_62_n3, CO => 
                           intadd_62_n2, S => intadd_62_SUM_1_port);
   intadd_62_U2 : FA_X1 port map( A => intadd_62_A_2_port, B => 
                           intadd_62_B_2_port, CI => intadd_62_n2, CO => 
                           intadd_62_n1, S => intadd_62_SUM_2_port);
   R_1302 : DFF_X2 port map( D => FP_B(1), CK => clk, Q => n10948, QN => n14594
                           );
   R_1465 : DFF_X1 port map( D => FP_A(11), CK => clk, Q => n8340, QN => n10689
                           );
   R_1324 : DFF_X1 port map( D => FP_A(1), CK => clk, Q => n14723, QN => n14586
                           );
   R_1566 : DFF_X1 port map( D => FP_A(5), CK => clk, Q => n14721, QN => n10882
                           );
   R_1455 : DFF_X1 port map( D => FP_A(15), CK => clk, Q => n14712, QN => 
                           n10717);
   R_1486 : DFF_X1 port map( D => FP_A(13), CK => clk, Q => n14463, QN => 
                           n10877);
   R_1482 : DFF_X1 port map( D => FP_A(3), CK => clk, Q => n_1075, QN => n10873
                           );
   R_1499 : DFF_X1 port map( D => FP_A(7), CK => clk, Q => n8355, QN => n10861)
                           ;
   I1_B_SIG_reg_2_inst : DFF_X1 port map( D => FP_B(2), CK => clk, Q => n14447,
                           QN => n381);
   R_1470 : DFF_X1 port map( D => FP_A(21), CK => clk, Q => n_1076, QN => 
                           n10879);
   R_1500 : DFF_X1 port map( D => n14710, CK => clk, Q => n14825, QN => n14507)
                           ;
   R_1494 : DFF_X1 port map( D => n14709, CK => clk, Q => n14759, QN => n_1077)
                           ;
   R_1280 : DFF_X1 port map( D => n14673, CK => clk, Q => n14715, QN => n_1078)
                           ;
   R_1350 : DFF_X1 port map( D => n14708, CK => clk, Q => n14760, QN => n_1079)
                           ;
   R_48 : DFF_X1 port map( D => n14906, CK => clk, Q => n14707, QN => n_1080);
   R_49 : DFF_X1 port map( D => n14904, CK => clk, Q => n14706, QN => n_1081);
   R_52 : DFF_X1 port map( D => n14886, CK => clk, Q => n14705, QN => n_1082);
   R_53 : DFF_X1 port map( D => n14887, CK => clk, Q => n14704, QN => n_1083);
   R_1517 : DFF_X1 port map( D => n14703, CK => clk, Q => n14789, QN => n_1084)
                           ;
   R_1224 : DFF_X1 port map( D => n10927, CK => clk, Q => SIG_in_27_port, QN =>
                           n10975);
   R_1258 : DFF_X1 port map( D => n10927, CK => clk, Q => n14730, QN => n_1085)
                           ;
   R_88 : DFF_X1 port map( D => n14701, CK => clk, Q => n14778, QN => n14499);
   R_95 : DFF_X1 port map( D => n14666, CK => clk, Q => n_1086, QN => n10716);
   R_107 : DFF_X1 port map( D => n14912, CK => clk, Q => n14700, QN => n_1087);
   R_120 : DFF_X1 port map( D => n14699, CK => clk, Q => n14735, QN => n10922);
   R_122 : DFF_X1 port map( D => n14698, CK => clk, Q => n14787, QN => n10682);
   R_1219 : DFF_X1 port map( D => n14697, CK => clk, Q => n14891, QN => n_1088)
                           ;
   R_153 : DFF_X1 port map( D => n14889, CK => clk, Q => n14696, QN => n_1089);
   R_154 : DFF_X1 port map( D => n14888, CK => clk, Q => n14695, QN => n_1090);
   R_212 : DFF_X1 port map( D => n14885, CK => clk, Q => n14694, QN => n_1091);
   R_227 : DFF_X1 port map( D => n14915, CK => clk, Q => n14693, QN => n_1092);
   R_229 : DFF_X1 port map( D => n14913, CK => clk, Q => n14692, QN => n_1093);
   R_236 : DFF_X1 port map( D => n14911, CK => clk, Q => n14691, QN => n_1094);
   R_256 : DFF_X1 port map( D => n14918, CK => clk, Q => n14690, QN => n_1095);
   R_269 : DFF_X1 port map( D => n14884, CK => clk, Q => n14689, QN => n_1096);
   R_286 : DFF_X1 port map( D => n14907, CK => clk, Q => n14688, QN => n_1097);
   R_315 : DFF_X1 port map( D => n2589, CK => clk, Q => n14687, QN => n_1098);
   R_316 : DFF_X1 port map( D => n8375, CK => clk, Q => n14686, QN => n_1099);
   R_317 : DFF_X1 port map( D => n10975, CK => clk, Q => n14685, QN => n_1100);
   R_326 : DFF_X1 port map( D => n14917, CK => clk, Q => n14684, QN => n_1101);
   R_339 : DFF_X1 port map( D => n14879, CK => clk, Q => n14683, QN => n_1102);
   R_437 : DFF_X1 port map( D => n14902, CK => clk, Q => n14682, QN => n_1103);
   R_666 : DFF_X1 port map( D => n14899, CK => clk, Q => n_1104, QN => n10808);
   R_686 : DFF_X1 port map( D => n14921, CK => clk, Q => n14681, QN => n_1105);
   R_801 : DFF_X1 port map( D => n2587, CK => clk, Q => n14680, QN => n_1106);
   R_832 : DFF_X1 port map( D => n14900, CK => clk, Q => n14679, QN => n14944);
   R_844 : DFF_X1 port map( D => n14898, CK => clk, Q => n14678, QN => n_1107);
   R_875 : DFF_X1 port map( D => n14446, CK => clk, Q => n14677, QN => n_1108);
   R_876 : DFF_X1 port map( D => n14920, CK => clk, Q => n14676, QN => n_1109);
   R_910 : DFF_X1 port map( D => n14446, CK => clk, Q => n14675, QN => n_1110);
   R_911 : DFF_X1 port map( D => n14920, CK => clk, Q => n14674, QN => n_1111);
   R_1521 : DFF_X1 port map( D => n14669, CK => clk, Q => n14740, QN => n14479)
                           ;
   R_1268 : DFF_X1 port map( D => n14668, CK => clk, Q => n14832, QN => n14492)
                           ;
   R_949 : DFF_X1 port map( D => n11430, CK => clk, Q => n14665, QN => n_1112);
   R_950 : DFF_X1 port map( D => n14920, CK => clk, Q => n14664, QN => n_1113);
   R_973 : DFF_X1 port map( D => FP_A(14), CK => clk, Q => n14734, QN => n_1114
                           );
   R_1574 : DFF_X1 port map( D => n384, CK => clk, Q => n14713, QN => n_1115);
   R_991 : DFF_X1 port map( D => n14847, CK => clk, Q => n14659, QN => n_1116);
   R_1421 : DFF_X1 port map( D => n14523, CK => clk, Q => n14770, QN => n14510)
                           ;
   R_1021 : DFF_X1 port map( D => n14817, CK => clk, Q => n14657, QN => n_1117)
                           ;
   R_1028 : DFF_X1 port map( D => n14862, CK => clk, Q => n14656, QN => n_1118)
                           ;
   R_1033 : DFF_X1 port map( D => n14808, CK => clk, Q => n14655, QN => n_1119)
                           ;
   R_1055 : DFF_X1 port map( D => n14652, CK => clk, Q => n14882, QN => n14480)
                           ;
   R_1059 : DFF_X1 port map( D => n14830, CK => clk, Q => n14651, QN => n_1120)
                           ;
   R_1061 : DFF_X1 port map( D => n14850, CK => clk, Q => n14650, QN => n_1121)
                           ;
   R_1063 : DFF_X1 port map( D => intadd_46_B_4_port, CK => clk, Q => n14649, 
                           QN => n14940);
   R_1064 : DFF_X1 port map( D => intadd_46_n2, CK => clk, Q => n14648, QN => 
                           n14941);
   R_1070 : DFF_X1 port map( D => n14865, CK => clk, Q => n14647, QN => n_1122)
                           ;
   R_1080 : DFF_X1 port map( D => I1_I1_N13, CK => clk, Q => n14881, QN => 
                           n14942);
   R_1084 : DFF_X1 port map( D => n14826, CK => clk, Q => n14645, QN => n_1123)
                           ;
   R_1090 : DFF_X1 port map( D => n14799, CK => clk, Q => n14644, QN => n_1124)
                           ;
   R_1104 : DFF_X1 port map( D => n14925, CK => clk, Q => n14643, QN => n_1125)
                           ;
   R_1106 : DFF_X1 port map( D => n14923, CK => clk, Q => n14642, QN => n_1126)
                           ;
   R_1112 : DFF_X1 port map( D => n14932, CK => clk, Q => n14641, QN => n_1127)
                           ;
   R_1115 : DFF_X1 port map( D => n14640, CK => clk, Q => n14840, QN => n14481)
                           ;
   R_1116 : DFF_X1 port map( D => n14639, CK => clk, Q => n14783, QN => n_1128)
                           ;
   R_1220 : DFF_X1 port map( D => n14491, CK => clk, Q => n14890, QN => n_1129)
                           ;
   R_1141 : DFF_X1 port map( D => n14790, CK => clk, Q => n14638, QN => n_1130)
                           ;
   R_1151 : DFF_X1 port map( D => n14836, CK => clk, Q => n14637, QN => n_1131)
                           ;
   R_1152 : DFF_X1 port map( D => n14835, CK => clk, Q => n14636, QN => n_1132)
                           ;
   R_1163 : DFF_X1 port map( D => intadd_66_n1, CK => clk, Q => n14635, QN => 
                           n_1133);
   R_1171 : DFF_X1 port map( D => n14797, CK => clk, Q => n14634, QN => n_1134)
                           ;
   R_1173 : DFF_X1 port map( D => n14810, CK => clk, Q => n14633, QN => n_1135)
                           ;
   R_1174 : DFF_X1 port map( D => n14809, CK => clk, Q => n14632, QN => n_1136)
                           ;
   R_1176 : DFF_X1 port map( D => n14828, CK => clk, Q => n14631, QN => n_1137)
                           ;
   R_1178 : DFF_X1 port map( D => n14774, CK => clk, Q => n14629, QN => n_1138)
                           ;
   R_1179 : DFF_X1 port map( D => n14773, CK => clk, Q => n14628, QN => n_1139)
                           ;
   R_1177 : DFF_X1 port map( D => n14775, CK => clk, Q => n14630, QN => n_1140)
                           ;
   R_1186 : DFF_X1 port map( D => n14834, CK => clk, Q => n14627, QN => n_1141)
                           ;
   R_1191 : DFF_X1 port map( D => n14860, CK => clk, Q => n14626, QN => n_1142)
                           ;
   R_1200 : DFF_X1 port map( D => n10676, CK => clk, Q => n14625, QN => n_1143)
                           ;
   R_1203 : DFF_X1 port map( D => n14875, CK => clk, Q => n14624, QN => n_1144)
                           ;
   R_1208 : DFF_X1 port map( D => intadd_61_n2, CK => clk, Q => n14623, QN => 
                           n_1145);
   R_1209 : DFF_X1 port map( D => intadd_61_n7, CK => clk, Q => n14622, QN => 
                           n_1146);
   R_1214 : DFF_X1 port map( D => n14838, CK => clk, Q => n14621, QN => n_1147)
                           ;
   R_1215 : DFF_X1 port map( D => n14837, CK => clk, Q => n14620, QN => n_1148)
                           ;
   R_1223 : DFF_X1 port map( D => n14873, CK => clk, Q => n14618, QN => n_1149)
                           ;
   R_1334 : DFF_X1 port map( D => n10927, CK => clk, Q => n14729, QN => n_1150)
                           ;
   R_1232 : DFF_X1 port map( D => n14746, CK => clk, Q => n14616, QN => n_1151)
                           ;
   R_1233 : DFF_X1 port map( D => n14745, CK => clk, Q => n14615, QN => n_1152)
                           ;
   R_1231 : DFF_X1 port map( D => n14747, CK => clk, Q => n14617, QN => n_1153)
                           ;
   R_1238 : DFF_X1 port map( D => n14857, CK => clk, Q => n14614, QN => n_1154)
                           ;
   R_1239 : DFF_X1 port map( D => n14870, CK => clk, Q => n14613, QN => n_1155)
                           ;
   R_1240 : DFF_X1 port map( D => n14856, CK => clk, Q => n14612, QN => n_1156)
                           ;
   R_1241 : DFF_X1 port map( D => n14855, CK => clk, Q => n14611, QN => n_1157)
                           ;
   R_1243 : DFF_X1 port map( D => n14767, CK => clk, Q => n14610, QN => n_1158)
                           ;
   R_1245 : DFF_X1 port map( D => n14919, CK => clk, Q => n14609, QN => n10929)
                           ;
   R_1120 : DFF_X1 port map( D => n10825, CK => clk, Q => n_1159, QN => n10826)
                           ;
   R_1249 : DFF_X1 port map( D => n14877, CK => clk, Q => n14608, QN => n_1160)
                           ;
   R_1259 : DFF_X1 port map( D => n14607, CK => clk, Q => n14895, QN => n_1161)
                           ;
   R_1545 : DFF_X1 port map( D => FP_A(3), CK => clk, Q => n14720, QN => n_1162
                           );
   R_1270 : DFF_X1 port map( D => n14604, CK => clk, Q => n14833, QN => n_1163)
                           ;
   R_1277 : DFF_X1 port map( D => n14732, CK => clk, Q => n14841, QN => n14460)
                           ;
   R_1281 : DFF_X1 port map( D => n14600, CK => clk, Q => n14878, QN => n_1164)
                           ;
   R_1283 : DFF_X1 port map( D => n14793, CK => clk, Q => n14599, QN => n_1165)
                           ;
   R_1290 : DFF_X1 port map( D => n14524, CK => clk, Q => n14781, QN => n_1166)
                           ;
   R_1303 : DFF_X1 port map( D => FP_B(1), CK => clk, Q => n14777, QN => n_1167
                           );
   R_1305 : DFF_X1 port map( D => FP_B(3), CK => clk, Q => n14785, QN => n_1168
                           );
   R_1310 : DFF_X1 port map( D => n14592, CK => clk, Q => n14737, QN => n_1169)
                           ;
   R_1311 : DFF_X1 port map( D => n14591, CK => clk, Q => n14819, QN => n_1170)
                           ;
   R_1308 : DFF_X1 port map( D => n14603, CK => clk, Q => n14456, QN => n14484)
                           ;
   R_1314 : DFF_X1 port map( D => n11676, CK => clk, Q => n14590, QN => n_1171)
                           ;
   R_1315 : DFF_X1 port map( D => n14852, CK => clk, Q => n14589, QN => n_1172)
                           ;
   R_1317 : DFF_X1 port map( D => n14843, CK => clk, Q => n14588, QN => n_1173)
                           ;
   R_1478 : DFF_X1 port map( D => FP_A(1), CK => clk, Q => n14784, QN => n_1174
                           );
   R_1322 : DFF_X1 port map( D => n14844, CK => clk, Q => n14587, QN => n_1175)
                           ;
   R_1325 : DFF_X1 port map( D => n14585, CK => clk, Q => n14771, QN => n14468)
                           ;
   R_1330 : DFF_X1 port map( D => n14582, CK => clk, Q => n14739, QN => n_1176)
                           ;
   R_1329 : DFF_X1 port map( D => n14583, CK => clk, Q => n14716, QN => n_1177)
                           ;
   R_1335 : DFF_X1 port map( D => n14581, CK => clk, Q => n14896, QN => n14495)
                           ;
   R_1337 : DFF_X1 port map( D => n14579, CK => clk, Q => n14741, QN => n_1178)
                           ;
   R_1338 : DFF_X1 port map( D => n14766, CK => clk, Q => n14578, QN => n_1179)
                           ;
   R_1339 : DFF_X1 port map( D => n14765, CK => clk, Q => n14577, QN => n_1180)
                           ;
   R_1340 : DFF_X1 port map( D => EXP_out_round_4_port, CK => clk, Q => n14576,
                           QN => n_1181);
   R_1341 : DFF_X1 port map( D => n14929, CK => clk, Q => n14575, QN => n_1182)
                           ;
   R_1343 : DFF_X1 port map( D => n14928, CK => clk, Q => n14574, QN => n_1183)
                           ;
   R_1349 : DFF_X1 port map( D => n14572, CK => clk, Q => n14738, QN => n_1184)
                           ;
   R_1355 : DFF_X1 port map( D => n14795, CK => clk, Q => n14570, QN => n_1185)
                           ;
   R_1358 : DFF_X1 port map( D => n14742, CK => clk, Q => n14568, QN => n_1186)
                           ;
   R_1361 : DFF_X1 port map( D => EXP_out_round_1_port, CK => clk, Q => n14566,
                           QN => n_1187);
   R_1363 : DFF_X1 port map( D => n14926, CK => clk, Q => n14565, QN => n_1188)
                           ;
   R_1360 : DFF_X1 port map( D => n14924, CK => clk, Q => n14567, QN => n_1189)
                           ;
   R_1364 : DFF_X1 port map( D => n14752, CK => clk, Q => n14564, QN => n_1190)
                           ;
   R_1365 : DFF_X1 port map( D => n14751, CK => clk, Q => n14563, QN => n_1191)
                           ;
   R_1367 : DFF_X1 port map( D => n14762, CK => clk, Q => n14562, QN => n_1192)
                           ;
   R_1422 : DFF_X1 port map( D => n14536, CK => clk, Q => n14880, QN => n14487)
                           ;
   R_1420 : DFF_X1 port map( D => I1_I0_N13, CK => clk, Q => n14718, QN => 
                           n14653);
   R_1221 : DFF_X1 port map( D => n14619, CK => clk, Q => n14894, QN => n_1193)
                           ;
   R_1495 : DFF_X2 port map( D => FP_B(0), CK => clk, Q => n14719, QN => n10864
                           );
   R_1546 : DFF_X2 port map( D => I1_I1_N13, CK => clk, Q => n14726, QN => 
                           n10841);
   R_1559 : DFF_X1 port map( D => FP_A(17), CK => clk, Q => n8353, QN => n10934
                           );
   R_1484 : DFF_X1 port map( D => FP_A(19), CK => clk, Q => n8339, QN => n10871
                           );
   R_1304 : DFF_X2 port map( D => FP_B(3), CK => clk, Q => n_1194, QN => n14593
                           );
   I1_B_EXP_reg_2_inst : DFF_X1 port map( D => FP_B(25), CK => clk, Q => 
                           B_EXP_2_port, QN => n14473);
   I1_A_EXP_reg_2_inst : DFF_X1 port map( D => FP_A(25), CK => clk, Q => 
                           A_EXP_2_port, QN => n14505);
   I3_EXP_out_round_reg_4_inst : DFF_X1 port map( D => I3_EXP_out_4_port, CK =>
                           clk, Q => EXP_out_round_4_port, QN => n14509);
   I3_EXP_out_round_reg_5_inst : DFF_X1 port map( D => I3_EXP_out_5_port, CK =>
                           clk, Q => n14498, QN => n8379);
   I2_SIG_in_reg_13_inst : DFF_X1 port map( D => I2_dtemp_33_port, CK => clk, Q
                           => n8345, QN => n14520);
   I2_SIG_in_reg_11_inst : DFF_X1 port map( D => I2_dtemp_31_port, CK => clk, Q
                           => n14512, QN => n8374);
   I2_SIG_in_reg_20_inst : DFF_X1 port map( D => n14938, CK => clk, Q => n14514
                           , QN => n2594);
   I2_SIG_in_reg_16_inst : DFF_X1 port map( D => n8409, CK => clk, Q => n14513,
                           QN => n2598);
   I2_SIG_in_reg_22_inst : DFF_X1 port map( D => I2_dtemp_42_port, CK => clk, Q
                           => n14516, QN => n2592);
   I2_SIG_in_reg_23_inst : DFF_X1 port map( D => I2_dtemp_43_port, CK => clk, Q
                           => n8347, QN => n14521);
   I2_SIG_in_reg_25_inst : DFF_X1 port map( D => n14935, CK => clk, Q => n14470
                           , QN => n2589);
   I2_SIG_in_reg_26_inst : DFF_X1 port map( D => n14916, CK => clk, Q => n8375,
                           QN => n14500);
   I2_SIG_in_reg_18_inst : DFF_X1 port map( D => n14934, CK => clk, Q => n14515
                           , QN => n2596);
   I1_B_SIG_reg_22_inst : DFF_X1 port map( D => FP_B(22), CK => clk, Q => n8331
                           , QN => n14459);
   R_1480 : DFF_X1 port map( D => FP_B(6), CK => clk, Q => n8352, QN => n10722)
                           ;
   R_945 : DFF_X1 port map( D => n14666, CK => clk, Q => n14727, QN => n_1195);
   R_935 : DFF_X1 port map( D => n14670, CK => clk, Q => n14780, QN => n10718);
   R_1435 : DFF_X1 port map( D => n14764, CK => clk, Q => n14526, QN => n_1196)
                           ;
   R_1434 : DFF_X1 port map( D => n14763, CK => clk, Q => n14527, QN => n_1197)
                           ;
   R_1433 : DFF_X1 port map( D => n14748, CK => clk, Q => n14528, QN => n_1198)
                           ;
   R_1429 : DFF_X1 port map( D => n14829, CK => clk, Q => n14529, QN => n_1199)
                           ;
   R_1428 : DFF_X1 port map( D => n14827, CK => clk, Q => n14530, QN => n_1200)
                           ;
   R_1427 : DFF_X1 port map( D => intadd_61_n6, CK => clk, Q => n14531, QN => 
                           n_1201);
   R_1426 : DFF_X1 port map( D => intadd_61_n1, CK => clk, Q => n14532, QN => 
                           n_1202);
   R_1425 : DFF_X1 port map( D => intadd_61_n5, CK => clk, Q => n14533, QN => 
                           n_1203);
   R_1424 : DFF_X1 port map( D => n14814, CK => clk, Q => n14534, QN => n_1204)
                           ;
   R_1423 : DFF_X1 port map( D => n14815, CK => clk, Q => n14535, QN => n_1205)
                           ;
   R_1419 : DFF_X1 port map( D => n14663, CK => clk, Q => n14883, QN => n_1206)
                           ;
   R_1418 : DFF_X1 port map( D => n14848, CK => clk, Q => n14537, QN => n_1207)
                           ;
   R_1416 : DFF_X1 port map( D => n14853, CK => clk, Q => n14538, QN => n_1208)
                           ;
   R_1415 : DFF_X1 port map( D => n14851, CK => clk, Q => n14539, QN => n_1209)
                           ;
   R_1412 : DFF_X1 port map( D => intadd_42_n11, CK => clk, Q => n14542, QN => 
                           n_1210);
   R_1411 : DFF_X1 port map( D => intadd_42_B_3_port, CK => clk, Q => n14543, 
                           QN => n_1211);
   R_1410 : DFF_X1 port map( D => intadd_42_A_3_port, CK => clk, Q => n14544, 
                           QN => n_1212);
   R_1409 : DFF_X1 port map( D => n14545, CK => clk, Q => n14893, QN => n_1213)
                           ;
   R_1408 : DFF_X1 port map( D => n14658, CK => clk, Q => n14892, QN => n_1214)
                           ;
   R_1407 : DFF_X1 port map( D => n14871, CK => clk, Q => n14546, QN => n_1215)
                           ;
   R_1405 : DFF_X1 port map( D => n14824, CK => clk, Q => n14547, QN => n_1216)
                           ;
   R_1404 : DFF_X1 port map( D => n14820, CK => clk, Q => n14548, QN => n_1217)
                           ;
   R_1399 : DFF_X1 port map( D => n14807, CK => clk, Q => n14550, QN => n_1218)
                           ;
   R_1398 : DFF_X1 port map( D => n14874, CK => clk, Q => n14551, QN => n_1219)
                           ;
   R_1396 : DFF_X1 port map( D => n14733, CK => clk, Q => n14736, QN => n_1220)
                           ;
   R_1492 : DFF_X1 port map( D => FP_A(8), CK => clk, Q => A_SIG_8_port, QN => 
                           n_1221);
   R_1510 : DFF_X1 port map( D => FP_A(7), CK => clk, Q => n14717, QN => n_1222
                           );
   R_1393 : DFF_X1 port map( D => n14867, CK => clk, Q => n14552, QN => n_1223)
                           ;
   R_1391 : DFF_X1 port map( D => n14903, CK => clk, Q => n14553, QN => n_1224)
                           ;
   R_1385 : DFF_X1 port map( D => n14846, CK => clk, Q => n14554, QN => n_1225)
                           ;
   R_1380 : DFF_X1 port map( D => n14858, CK => clk, Q => n14555, QN => n_1226)
                           ;
   R_1379 : DFF_X1 port map( D => n14859, CK => clk, Q => n14556, QN => n_1227)
                           ;
   R_1378 : DFF_X1 port map( D => n14557, CK => clk, Q => n14788, QN => n10973)
                           ;
   R_1376 : DFF_X1 port map( D => n14822, CK => clk, Q => n14558, QN => n_1228)
                           ;
   R_1372 : DFF_X1 port map( D => n14821, CK => clk, Q => n14559, QN => n_1229)
                           ;
   R_1370 : DFF_X1 port map( D => n14816, CK => clk, Q => n14560, QN => n_1230)
                           ;
   R_1368 : DFF_X1 port map( D => n14761, CK => clk, Q => n14561, QN => n_1231)
                           ;
   R_1491 : DFF_X1 port map( D => FP_A(9), CK => clk, Q => n8338, QN => n10866)
                           ;
   R_1352 : DFF_X2 port map( D => n14571, CK => clk, Q => n14813, QN => n14483)
                           ;
   R_1347 : DFF_X1 port map( D => FP_B(12), CK => clk, Q => n4381, QN => n14455
                           );
   R_929 : DFF_X2 port map( D => n14672, CK => clk, Q => n14779, QN => n10733);
   R_1454 : DFF_X1 port map( D => FP_B(18), CK => clk, Q => n12125, QN => 
                           n_1232);
   R_1458 : DFF_X1 port map( D => n10883, CK => clk, Q => n12639, QN => n10637)
                           ;
   R_1462 : DFF_X1 port map( D => n10881, CK => clk, Q => n11097, QN => n_1233)
                           ;
   R_1464 : DFF_X1 port map( D => FP_A(9), CK => clk, Q => n12124, QN => n_1234
                           );
   R_1469 : DFF_X1 port map( D => n10880, CK => clk, Q => n13362, QN => n10630)
                           ;
   R_1474 : DFF_X1 port map( D => n10876, CK => clk, Q => n11164, QN => n_1235)
                           ;
   R_1475 : DFF_X1 port map( D => n14580, CK => clk, Q => n11861, QN => n_1236)
                           ;
   R_1476 : DFF_X1 port map( D => n10875, CK => clk, Q => n10983, QN => n_1237)
                           ;
   R_1481 : DFF_X1 port map( D => FP_B(6), CK => clk, Q => n13924, QN => n_1238
                           );
   R_1483 : DFF_X1 port map( D => n10872, CK => clk, Q => n13967, QN => n10634)
                           ;
   R_1485 : DFF_X1 port map( D => n10870, CK => clk, Q => n11283, QN => n_1239)
                           ;
   R_1488 : DFF_X1 port map( D => n10868, CK => clk, Q => n12173, QN => n_1240)
                           ;
   R_1490 : DFF_X1 port map( D => n13528, CK => clk, Q => n10867, QN => n_1241)
                           ;
   R_1493 : DFF_X1 port map( D => n10865, CK => clk, Q => n11385, QN => n10640)
                           ;
   R_1496 : DFF_X1 port map( D => n10863, CK => clk, Q => n11305, QN => n_1242)
                           ;
   R_1498 : DFF_X1 port map( D => n10862, CK => clk, Q => n_1243, QN => n10714)
                           ;
   R_1501 : DFF_X1 port map( D => n10860, CK => clk, Q => n11149, QN => n10642)
                           ;
   R_1502 : DFF_X1 port map( D => n13574, CK => clk, Q => n10859, QN => n_1244)
                           ;
   R_1503 : DFF_X1 port map( D => n14187, CK => clk, Q => n10858, QN => n_1245)
                           ;
   R_1511 : DFF_X1 port map( D => n10856, CK => clk, Q => n11043, QN => n10638)
                           ;
   R_1512 : DFF_X1 port map( D => n13578, CK => clk, Q => n10855, QN => n_1246)
                           ;
   R_1513 : DFF_X1 port map( D => n13577, CK => clk, Q => n10854, QN => n_1247)
                           ;
   R_1516 : DFF_X1 port map( D => n10852, CK => clk, Q => n11369, QN => n_1248)
                           ;
   R_1518 : DFF_X1 port map( D => n10851, CK => clk, Q => n10952, QN => n_1249)
                           ;
   R_1524 : DFF_X1 port map( D => FP_B(11), CK => clk, Q => n13273, QN => 
                           n_1250);
   R_1525 : DFF_X1 port map( D => n13527, CK => clk, Q => n10849, QN => n_1251)
                           ;
   R_1526 : DFF_X1 port map( D => n13526, CK => clk, Q => n10848, QN => n_1252)
                           ;
   R_1527 : DFF_X1 port map( D => n14431, CK => clk, Q => n10847, QN => n_1253)
                           ;
   R_1529 : DFF_X1 port map( D => n14430, CK => clk, Q => n10846, QN => n_1254)
                           ;
   R_1532 : DFF_X1 port map( D => n11827, CK => clk, Q => n10845, QN => n_1255)
                           ;
   R_1534 : DFF_X1 port map( D => n14102, CK => clk, Q => n10844, QN => n_1256)
                           ;
   R_1535 : DFF_X1 port map( D => n14101, CK => clk, Q => n10843, QN => n_1257)
                           ;
   R_1538 : DFF_X1 port map( D => n10842, CK => clk, Q => n_1258, QN => n10631)
                           ;
   R_1540 : DFF_X1 port map( D => FP_B(7), CK => clk, Q => n10905, QN => n_1259
                           );
   R_1542 : DFF_X1 port map( D => FP_B(9), CK => clk, Q => n11738, QN => n_1260
                           );
   R_1547 : DFF_X1 port map( D => n10840, CK => clk, Q => n12023, QN => n_1261)
                           ;
   R_1548 : DFF_X1 port map( D => n13217, CK => clk, Q => n10839, QN => n_1262)
                           ;
   R_1549 : DFF_X1 port map( D => n13218, CK => clk, Q => n10838, QN => n_1263)
                           ;
   R_1551 : DFF_X1 port map( D => n14435, CK => clk, Q => n10837, QN => n_1264)
                           ;
   R_1552 : DFF_X1 port map( D => n14434, CK => clk, Q => n10836, QN => n_1265)
                           ;
   R_1554 : DFF_X1 port map( D => n10835, CK => clk, Q => n_1266, QN => n10635)
                           ;
   R_1560 : DFF_X1 port map( D => n10834, CK => clk, Q => n11225, QN => n10636)
                           ;
   R_1562 : DFF_X1 port map( D => n14441, CK => clk, Q => n10833, QN => n_1267)
                           ;
   R_1563 : DFF_X1 port map( D => n14440, CK => clk, Q => n10832, QN => n_1268)
                           ;
   R_1568 : DFF_X1 port map( D => n10830, CK => clk, Q => n11488, QN => n_1269)
                           ;
   R_1569 : DFF_X1 port map( D => FP_A(5), CK => clk, Q => n11487, QN => n_1270
                           );
   R_1571 : DFF_X1 port map( D => n10705, CK => clk, Q => n10829, QN => n_1271)
                           ;
   R_1572 : DFF_X1 port map( D => n13627, CK => clk, Q => n10828, QN => n_1272)
                           ;
   R_1573 : DFF_X1 port map( D => n13626, CK => clk, Q => n10827, QN => n_1273)
                           ;
   R_1575 : DFF_X1 port map( D => n384, CK => clk, Q => n12671, QN => n_1274);
   R_1592 : DFF_X1 port map( D => intadd_63_SUM_2_port, CK => clk, Q => n10824,
                           QN => n_1275);
   R_1593 : DFF_X1 port map( D => intadd_46_SUM_3_port, CK => clk, Q => n10823,
                           QN => n_1276);
   R_1594 : DFF_X1 port map( D => intadd_62_n1, CK => clk, Q => n10822, QN => 
                           n10821);
   R_1595 : DFF_X1 port map( D => intadd_46_SUM_2_port, CK => clk, Q => n10820,
                           QN => n_1277);
   R_1596 : DFF_X1 port map( D => intadd_62_SUM_2_port, CK => clk, Q => n10819,
                           QN => n_1278);
   R_1597 : DFF_X1 port map( D => n14905, CK => clk, Q => n10818, QN => n_1279)
                           ;
   R_1598 : DFF_X1 port map( D => n14897, CK => clk, Q => n10817, QN => n_1280)
                           ;
   R_1599 : DFF_X1 port map( D => n14757, CK => clk, Q => n10816, QN => n10643)
                           ;
   R_1600 : DFF_X1 port map( D => n14758, CK => clk, Q => n10815, QN => n10632)
                           ;
   R_1602 : DFF_X1 port map( D => intadd_66_SUM_2_port, CK => clk, Q => n10814,
                           QN => n_1281);
   R_1603 : DFF_X1 port map( D => n13214, CK => clk, Q => n10813, QN => n_1282)
                           ;
   R_1604 : DFF_X1 port map( D => n10937, CK => clk, Q => n10812, QN => n_1283)
                           ;
   R_1605 : DFF_X1 port map( D => n14525, CK => clk, Q => n10811, QN => n14943)
                           ;
   R_1606 : DFF_X1 port map( D => n2567, CK => clk, Q => n10807, QN => n10806);
   R_1607 : DFF_X1 port map( D => n2565, CK => clk, Q => n10805, QN => n_1284);
   R_1608 : DFF_X1 port map( D => n2556, CK => clk, Q => n10804, QN => n_1285);
   R_1609 : DFF_X1 port map( D => n2568, CK => clk, Q => n10803, QN => n_1286);
   R_1610 : DFF_X1 port map( D => n2557, CK => clk, Q => n10802, QN => n_1287);
   R_1611 : DFF_X1 port map( D => n2569, CK => clk, Q => n10801, QN => n_1288);
   R_1612 : DFF_X1 port map( D => n2558, CK => clk, Q => n10800, QN => n_1289);
   R_1613 : DFF_X1 port map( D => n2570, CK => clk, Q => n10799, QN => n_1290);
   R_1614 : DFF_X1 port map( D => n2559, CK => clk, Q => n10798, QN => n_1291);
   R_1615 : DFF_X1 port map( D => n2571, CK => clk, Q => n10797, QN => n_1292);
   R_1616 : DFF_X1 port map( D => n2560, CK => clk, Q => n10796, QN => n_1293);
   R_1617 : DFF_X1 port map( D => n2572, CK => clk, Q => n10795, QN => n_1294);
   R_1618 : DFF_X1 port map( D => n2561, CK => clk, Q => n10794, QN => n_1295);
   R_1619 : DFF_X1 port map( D => n2573, CK => clk, Q => n10793, QN => n_1296);
   R_1620 : DFF_X1 port map( D => n2562, CK => clk, Q => n10792, QN => n_1297);
   R_1621 : DFF_X1 port map( D => n2574, CK => clk, Q => n10791, QN => n_1298);
   R_1622 : DFF_X1 port map( D => n2563, CK => clk, Q => n10790, QN => n_1299);
   R_1623 : DFF_X1 port map( D => n14910, CK => clk, Q => n10789, QN => n_1300)
                           ;
   R_1624 : DFF_X1 port map( D => n14908, CK => clk, Q => n10788, QN => n_1301)
                           ;
   R_1625 : DFF_X1 port map( D => n14901, CK => clk, Q => n10787, QN => n_1302)
                           ;
   R_1626 : DFF_X1 port map( D => n14876, CK => clk, Q => n10786, QN => n_1303)
                           ;
   R_1627 : DFF_X1 port map( D => n14864, CK => clk, Q => n10785, QN => n_1304)
                           ;
   R_1628 : DFF_X1 port map( D => n14866, CK => clk, Q => n10784, QN => n_1305)
                           ;
   R_1629 : DFF_X1 port map( D => n14872, CK => clk, Q => n10783, QN => n_1306)
                           ;
   R_1630 : DFF_X1 port map( D => n14854, CK => clk, Q => n10782, QN => n_1307)
                           ;
   R_1631 : DFF_X1 port map( D => n14849, CK => clk, Q => n10781, QN => n_1308)
                           ;
   R_1632 : DFF_X1 port map( D => n14812, CK => clk, Q => n10780, QN => n_1309)
                           ;
   R_1633 : DFF_X1 port map( D => n14806, CK => clk, Q => n10779, QN => n_1310)
                           ;
   R_1634 : DFF_X1 port map( D => n14798, CK => clk, Q => n10778, QN => n_1311)
                           ;
   R_1635 : DFF_X1 port map( D => n14800, CK => clk, Q => n10777, QN => n_1312)
                           ;
   R_1636 : DFF_X1 port map( D => n14754, CK => clk, Q => n10776, QN => n10775)
                           ;
   R_1637 : DFF_X1 port map( D => n14869, CK => clk, Q => n10774, QN => n10773)
                           ;
   R_1638 : DFF_X1 port map( D => n14863, CK => clk, Q => n10772, QN => n_1313)
                           ;
   R_1639 : DFF_X1 port map( D => n14868, CK => clk, Q => n10771, QN => n_1314)
                           ;
   R_1640 : DFF_X1 port map( D => n14839, CK => clk, Q => n10770, QN => n_1315)
                           ;
   R_1641 : DFF_X1 port map( D => n14845, CK => clk, Q => n10769, QN => n_1316)
                           ;
   R_1642 : DFF_X1 port map( D => n14802, CK => clk, Q => n10768, QN => n_1317)
                           ;
   R_1643 : DFF_X1 port map( D => n13601, CK => clk, Q => n10767, QN => n_1318)
                           ;
   R_1644 : DFF_X1 port map( D => n13602, CK => clk, Q => n10766, QN => n_1319)
                           ;
   R_1645 : DFF_X1 port map( D => n10686, CK => clk, Q => n10765, QN => n_1320)
                           ;
   R_1646 : DFF_X1 port map( D => n14803, CK => clk, Q => n10764, QN => n_1321)
                           ;
   R_1647 : DFF_X1 port map( D => n14486, CK => clk, Q => n10763, QN => n_1322)
                           ;
   R_1648 : DFF_X1 port map( D => n14485, CK => clk, Q => n10762, QN => n_1323)
                           ;
   R_1649 : DFF_X1 port map( D => n14462, CK => clk, Q => n10761, QN => n_1324)
                           ;
   R_1650 : DFF_X1 port map( D => n14461, CK => clk, Q => n10760, QN => n_1325)
                           ;
   R_1651 : DFF_X1 port map( D => n14914, CK => clk, Q => n10759, QN => n_1326)
                           ;
   R_1652 : DFF_X1 port map( D => n14909, CK => clk, Q => n10758, QN => n_1327)
                           ;
   R_1653 : DFF_X1 port map( D => n13603, CK => clk, Q => n10757, QN => n_1328)
                           ;
   R_1654 : DFF_X1 port map( D => n13616, CK => clk, Q => n10756, QN => n_1329)
                           ;
   R_1655 : DFF_X1 port map( D => n13618, CK => clk, Q => n10755, QN => n_1330)
                           ;
   R_1656 : DFF_X1 port map( D => n14861, CK => clk, Q => n10754, QN => n10753)
                           ;
   R_1657 : DFF_X1 port map( D => n14769, CK => clk, Q => n10752, QN => n10751)
                           ;
   R_1658 : DFF_X1 port map( D => n11483, CK => clk, Q => n10750, QN => n_1331)
                           ;
   R_1659 : DFF_X1 port map( D => n14801, CK => clk, Q => n10749, QN => n_1332)
                           ;
   R_1660 : DFF_X1 port map( D => n14755, CK => clk, Q => n10748, QN => n_1333)
                           ;
   R_1662 : DFF_X1 port map( D => n10970, CK => clk, Q => n10747, QN => n_1334)
                           ;
   R_1663 : DFF_X1 port map( D => n10936, CK => clk, Q => n10746, QN => n_1335)
                           ;
   I1_B_SIG_reg_13_inst : DFF_X1 port map( D => FP_B(13), CK => clk, Q => n8326
                           , QN => n14477);
   R_1289 : DFF_X1 port map( D => n14595, CK => clk, Q => n14818, QN => n10724)
                           ;
   R_1472 : DFF_X1 port map( D => FP_A(11), CK => clk, Q => n14725, QN => 
                           n10920);
   R_1414 : DFF_X2 port map( D => n14540, CK => clk, Q => n14728, QN => n_1336)
                           ;
   R_972 : DFF_X1 port map( D => n14660, CK => clk, Q => n10641, QN => n10704);
   R_1509 : DFF_X1 port map( D => n14662, CK => clk, Q => n14782, QN => n10857)
                           ;
   R_1514 : DFF_X1 port map( D => FP_B(5), CK => clk, Q => n14731, QN => n10950
                           );
   R_1345 : DFF_X1 port map( D => n10727, CK => clk, Q => n14573, QN => n_1337)
                           ;
   R_1309 : DFF_X2 port map( D => FP_B(8), CK => clk, Q => B_SIG_8_port, QN => 
                           n14469);
   R_1291 : DFF_X1 port map( D => FP_B(5), CK => clk, Q => n8401, QN => n14448)
                           ;
   R_1522 : DFF_X1 port map( D => n10850, CK => clk, Q => n14114, QN => n10633)
                           ;
   U3571 : AND2_X1 port map( A1 => n11780, A2 => n11779, ZN => n13618);
   U3572 : NAND2_X1 port map( A1 => n14201, A2 => n10721, ZN => n10618);
   U3573 : INV_X1 port map( A => n11668, ZN => n10620);
   U3574 : INV_X1 port map( A => n13507, ZN => n13504);
   U3575 : INV_X1 port map( A => n11621, ZN => n10608);
   U3576 : INV_X1 port map( A => n11622, ZN => n10609);
   U3577 : NAND2_X1 port map( A1 => n10601, A2 => n12627, ZN => n13097);
   U3578 : AND2_X1 port map( A1 => n11605, A2 => n14723, ZN => n11596);
   U3579 : NOR2_X1 port map( A1 => n13442, A2 => n14025, ZN => n10602);
   U3580 : XNOR2_X1 port map( A => n14717, B => n14469, ZN => n11152);
   U3581 : OR2_X1 port map( A1 => n14881, A2 => n14492, ZN => n10626);
   U3585 : NAND2_X1 port map( A1 => n12777, A2 => n12776, ZN => n12778);
   U3586 : AND2_X1 port map( A1 => n12807, A2 => n12806, ZN => n12808);
   U3587 : NAND2_X1 port map( A1 => n10609, A2 => n10608, ZN => n13507);
   U3588 : INV_X1 port map( A => n12778, ZN => n12815);
   U3592 : XNOR2_X1 port map( A => n11286, B => n10603, ZN => n10924);
   U3593 : NAND2_X1 port map( A1 => n10619, A2 => n10618, ZN => n13560);
   U3594 : AOI21_X1 port map( B1 => n12625, B2 => n13279, A => n10602, ZN => 
                           n10601);
   U3596 : XNOR2_X1 port map( A => n10662, B => n11073, ZN => n14062);
   U3598 : NOR2_X1 port map( A1 => n13598, A2 => n13520, ZN => n10615);
   U3601 : AOI22_X2 port map( A1 => n13378, A2 => n13416, B1 => n13376, B2 => 
                           n13377, ZN => n10670);
   U3603 : BUF_X2 port map( A => B_SIG_9_port, Z => n13368);
   U3604 : INV_X1 port map( A => n13493, ZN => n10603);
   U3605 : AND2_X2 port map( A1 => n11842, A2 => n11841, ZN => n12032);
   U3606 : NAND2_X2 port map( A1 => n12402, A2 => n12403, ZN => n12578);
   U3607 : AND2_X2 port map( A1 => n13440, A2 => n13439, ZN => n13677);
   U3608 : NAND2_X2 port map( A1 => n14778, A2 => n10873, ZN => n11201);
   U3611 : INV_X2 port map( A => n14469, ZN => n11703);
   U3613 : NOR2_X2 port map( A1 => n12550, A2 => n12557, ZN => n12519);
   U3614 : BUF_X1 port map( A => n11418, Z => n11900);
   U3615 : NAND2_X1 port map( A1 => n10597, A2 => n13540, ZN => n13543);
   U3616 : INV_X1 port map( A => n13539, ZN => n10597);
   U3617 : AND2_X2 port map( A1 => n13496, A2 => n13497, ZN => n13539);
   U3618 : AND2_X2 port map( A1 => n11405, A2 => n13885, ZN => n11555);
   U3619 : NOR2_X1 port map( A1 => n11274, A2 => n10604, ZN => n11282);
   U3620 : NAND2_X1 port map( A1 => n14841, A2 => n8339, ZN => n10737);
   U3621 : BUF_X1 port map( A => n11650, Z => n11651);
   U3623 : NOR2_X1 port map( A1 => n11322, A2 => n14740, ZN => n10598);
   U3624 : INV_X1 port map( A => n11634, ZN => n13050);
   U3625 : NAND2_X1 port map( A1 => n12152, A2 => n11634, ZN => n11637);
   U3627 : NAND2_X1 port map( A1 => n11631, A2 => n10971, ZN => n10599);
   U3628 : NAND2_X1 port map( A1 => n11632, A2 => n11633, ZN => n10600);
   U3629 : BUF_X2 port map( A => n10737, Z => n10736);
   U3630 : AND2_X2 port map( A1 => n10691, A2 => n13242, ZN => n13406);
   U3631 : NAND2_X1 port map( A1 => n10607, A2 => n10605, ZN => n10604);
   U3632 : NAND2_X1 port map( A1 => n12243, A2 => n14464, ZN => n10605);
   U3634 : NAND2_X1 port map( A1 => n11513, A2 => n11272, ZN => n10607);
   U3635 : NAND2_X1 port map( A1 => n10610, A2 => n12992, ZN => n12994);
   U3636 : NAND2_X1 port map( A1 => n12187, A2 => n12186, ZN => n10610);
   U3637 : NAND2_X1 port map( A1 => n10613, A2 => n10611, ZN => n11092);
   U3638 : NAND2_X1 port map( A1 => n14466, A2 => n14020, ZN => n10611);
   U3640 : NAND2_X1 port map( A1 => n10939, A2 => n13282, ZN => n10613);
   U3641 : OR2_X2 port map( A1 => n12253, A2 => n14895, ZN => n12252);
   U3642 : NOR2_X2 port map( A1 => n13265, A2 => n14483, ZN => n13323);
   U3643 : OAI21_X1 port map( B1 => n14965, B2 => n10615, A => n10614, ZN => 
                           n13549);
   U3644 : NAND2_X1 port map( A1 => n13520, A2 => n13598, ZN => n10614);
   U3646 : NAND2_X1 port map( A1 => n10617, A2 => n13879, ZN => n11384);
   U3647 : NAND2_X1 port map( A1 => n13878, A2 => n13877, ZN => n10617);
   U3648 : AND3_X2 port map( A1 => n14074, A2 => n13131, A3 => n13151, ZN => 
                           n14100);
   U3649 : AND2_X2 port map( A1 => n13109, A2 => n13111, ZN => n12922);
   U3650 : OAI21_X1 port map( B1 => n10721, B2 => n14201, A => n14207, ZN => 
                           n10619);
   U3651 : XNOR2_X1 port map( A => n11258, B => n10620, ZN => n10740);
   U3652 : NAND2_X1 port map( A1 => n10623, A2 => n10621, ZN => n11836);
   U3653 : NAND2_X1 port map( A1 => n11043, A2 => n14466, ZN => n10621);
   U3655 : NAND2_X1 port map( A1 => n11957, A2 => n13282, ZN => n10623);
   U3656 : XNOR2_X2 port map( A => n12269, B => n10777, ZN => n12322);
   U3658 : AOI22_X2 port map( A1 => n11459, A2 => n11718, B1 => n11458, B2 => 
                           n10741, ZN => n11476);
   U3660 : NAND2_X1 port map( A1 => n10624, A2 => n12787, ZN => n12790);
   U3661 : NAND2_X1 port map( A1 => n10958, A2 => n13295, ZN => n10624);
   U3663 : NAND2_X1 port map( A1 => n13449, A2 => n10626, ZN => n10625);
   U3664 : NOR2_X1 port map( A1 => n12783, A2 => n14942, ZN => n10627);
   U3665 : XNOR2_X1 port map( A => n13256, B => n12811, ZN => n10912);
   U3667 : AND2_X1 port map( A1 => n11645, A2 => n11644, ZN => n12156);
   U3668 : AOI22_X1 port map( A1 => n11107, A2 => n11550, B1 => n11106, B2 => 
                           n11105, ZN => n11549);
   U3669 : OR2_X1 port map( A1 => n12004, A2 => n12005, ZN => n12926);
   U3670 : NAND2_X1 port map( A1 => n13189, A2 => n13188, ZN => n13220);
   U3671 : OAI22_X1 port map( A1 => n10661, A2 => n11685, B1 => n11684, B2 => 
                           n14062, ZN => n11828);
   U3672 : AND2_X1 port map( A1 => n12131, A2 => n12130, ZN => n10644);
   U3673 : NOR2_X2 port map( A1 => n13968, A2 => n10634, ZN => n11096);
   U3674 : AND2_X2 port map( A1 => n11908, A2 => n11907, ZN => n12007);
   U3676 : CLKBUF_X1 port map( A => n11215, Z => n11216);
   U3677 : OR2_X1 port map( A1 => n13388, A2 => n10670, ZN => n10669);
   U3678 : AND2_X1 port map( A1 => n13433, A2 => n13429, ZN => n13436);
   U3680 : BUF_X1 port map( A => n8326, Z => n10743);
   U3681 : NAND2_X1 port map( A1 => n10857, A2 => n10861, ZN => n10680);
   U3682 : AND2_X2 port map( A1 => n8353, A2 => n10983, ZN => n12146);
   U3683 : BUF_X1 port map( A => n14466, Z => n10726);
   U3684 : BUF_X1 port map( A => n11097, Z => n13920);
   U3687 : BUF_X1 port map( A => n8333, Z => n13485);
   U3689 : CLKBUF_X2 port map( A => n8331, Z => n13261);
   U3690 : BUF_X2 port map( A => n14118, Z => n10645);
   U3691 : NAND2_X2 port map( A1 => n14759, A2 => n10871, ZN => n13442);
   U3692 : BUF_X2 port map( A => n11283, Z => n12163);
   U3693 : INV_X1 port map( A => FP_A(3), ZN => n14541);
   U3694 : INV_X1 port map( A => FP_A(10), ZN => n14667);
   U3695 : INV_X1 port map( A => FP_A(19), ZN => n14722);
   U3696 : INV_X1 port map( A => FP_A(21), ZN => n14673);
   U3697 : INV_X1 port map( A => FP_A(7), ZN => n14724);
   U3698 : INV_X1 port map( A => FP_A(13), ZN => n14580);
   U3699 : INV_X1 port map( A => FP_A(14), ZN => n14661);
   U3700 : INV_X1 port map( A => FP_A(5), ZN => n14596);
   U3701 : INV_X1 port map( A => FP_A(16), ZN => n14602);
   U3702 : INV_X1 port map( A => FP_A(9), ZN => n14605);
   U3703 : INV_X1 port map( A => FP_B(14), ZN => n359);
   U3704 : INV_X1 port map( A => FP_B(16), ZN => n360);
   U3705 : INV_X1 port map( A => FP_B(0), ZN => n2638);
   U3706 : OR2_X1 port map( A1 => n14811, A2 => n13551, ZN => n14094);
   U3707 : NAND2_X1 port map( A1 => n10650, A2 => n10649, ZN => intadd_46_n2);
   U3708 : AND2_X1 port map( A1 => n11808, A2 => n11807, ZN => n13616);
   U3710 : XNOR2_X1 port map( A => n10651, B => intadd_46_n3, ZN => 
                           intadd_46_SUM_3_port);
   U3711 : XOR2_X1 port map( A => n13832, B => n14291, Z => 
                           intadd_63_SUM_2_port);
   U3712 : OAI211_X1 port map( C1 => n14045, C2 => n14046, A => n14047, B => 
                           n10654, ZN => n14050);
   U3713 : NAND2_X1 port map( A1 => n10668, A2 => n10667, ZN => n13392);
   U3714 : AOI21_X1 port map( B1 => n13834, B2 => n13835, A => n13831, ZN => 
                           n14291);
   U3715 : INV_X1 port map( A => n12993, ZN => n10646);
   U3716 : XNOR2_X1 port map( A => n13636, B => n10674, ZN => n14258);
   U3717 : CLKBUF_X1 port map( A => n13187, Z => n13219);
   U3718 : CLKBUF_X1 port map( A => n13160, Z => n13161);
   U3719 : NAND2_X1 port map( A1 => n13387, A2 => n10669, ZN => n10668);
   U3720 : AND2_X1 port map( A1 => n11684, A2 => n14062, ZN => n10661);
   U3721 : XNOR2_X1 port map( A => n10672, B => n13670, ZN => n13671);
   U3722 : INV_X1 port map( A => n13437, ZN => n10674);
   U3723 : OAI21_X1 port map( B1 => n13436, B2 => n13430, A => n10675, ZN => 
                           n13437);
   U3724 : AOI22_X1 port map( A1 => n11509, A2 => n11542, B1 => n11540, B2 => 
                           n11541, ZN => n13162);
   U3725 : OR2_X1 port map( A1 => n13830, A2 => n13829, ZN => n13834);
   U3726 : OR2_X1 port map( A1 => n14049, A2 => n14048, ZN => n10654);
   U3727 : XNOR2_X1 port map( A => n13992, B => n13993, ZN => n14045);
   U3728 : OR2_X1 port map( A1 => n11327, A2 => n11328, ZN => n11563);
   U3730 : AND3_X1 port map( A1 => n13752, A2 => n14704, A3 => n14705, ZN => 
                           n10696);
   U3731 : XNOR2_X1 port map( A => n13227, B => n10658, ZN => n13394);
   U3732 : NAND2_X1 port map( A1 => n13435, A2 => n13434, ZN => n10675);
   U3733 : XNOR2_X1 port map( A => n11491, B => n10893, ZN => n11686);
   U3734 : INV_X1 port map( A => n11679, ZN => n10647);
   U3735 : XNOR2_X1 port map( A => n10671, B => n10720, ZN => n13670);
   U3736 : XNOR2_X1 port map( A => n12138, B => n10644, ZN => n13036);
   U3737 : AND2_X1 port map( A1 => n12439, A2 => n14683, ZN => n13752);
   U3738 : XNOR2_X1 port map( A => n10966, B => n11789, ZN => n11820);
   U3739 : XNOR2_X1 port map( A => n13415, B => n10673, ZN => n13669);
   U3740 : AOI22_X1 port map( A1 => n10657, A2 => n13009, B1 => n13007, B2 => 
                           n13008, ZN => n13138);
   U3741 : OAI21_X1 port map( B1 => n13508, B2 => n13507, A => n10903, ZN => 
                           n13639);
   U3742 : INV_X1 port map( A => n11252, ZN => n11251);
   U3743 : OR2_X1 port map( A1 => n11037, A2 => n11036, ZN => n12621);
   U3744 : XNOR2_X1 port map( A => n13414, B => n13411, ZN => n10671);
   U3745 : CLKBUF_X1 port map( A => n11405, Z => n13884);
   U3746 : INV_X1 port map( A => n12030, ZN => n10657);
   U3747 : OR2_X1 port map( A1 => n11130, A2 => n11129, ZN => n11136);
   U3748 : AND2_X1 port map( A1 => n13432, A2 => n13431, ZN => n13435);
   U3749 : INV_X1 port map( A => n10974, ZN => n10655);
   U3750 : OR2_X1 port map( A1 => n11100, A2 => n11099, ZN => n11553);
   U3751 : AND2_X1 port map( A1 => n12182, A2 => n10664, ZN => n12997);
   U3752 : OAI21_X1 port map( B1 => n10665, B2 => n11247, A => n11249, ZN => 
                           n11252);
   U3753 : XNOR2_X1 port map( A => n11259, B => n11261, ZN => n10652);
   U3754 : OAI21_X1 port map( B1 => n14121, B2 => n13444, A => n13443, ZN => 
                           n13651);
   U3756 : NOR2_X1 port map( A1 => n10985, A2 => n10984, ZN => n13072);
   U3757 : AND2_X1 port map( A1 => n10982, A2 => n10981, ZN => n13073);
   U3758 : NOR2_X1 port map( A1 => n12177, A2 => n12176, ZN => n12996);
   U3759 : OR2_X1 port map( A1 => n12028, A2 => n12029, ZN => n12030);
   U3760 : AND2_X1 port map( A1 => n11362, A2 => n13881, ZN => n10955);
   U3761 : NAND2_X1 port map( A1 => n11836, A2 => n11835, ZN => n12034);
   U3763 : OR2_X1 port map( A1 => n12148, A2 => n12147, ZN => n12149);
   U3764 : AND2_X1 port map( A1 => n12137, A2 => n12136, ZN => n12138);
   U3765 : NAND2_X1 port map( A1 => n11003, A2 => n12174, ZN => n11004);
   U3766 : INV_X1 port map( A => n13965, ZN => n13922);
   U3767 : OAI22_X1 port map( A1 => n11601, A2 => n14483, B1 => n11600, B2 => 
                           n11599, ZN => n10898);
   U3768 : NAND2_X1 port map( A1 => n11248, A2 => n10666, ZN => n10665);
   U3769 : NAND2_X1 port map( A1 => n13284, A2 => n12174, ZN => n13285);
   U3771 : BUF_X1 port map( A => n11201, Z => n13984);
   U3772 : INV_X1 port map( A => n10704, ZN => n10745);
   U3773 : AOI21_X1 port map( B1 => n11597, B2 => n10861, A => n12010, ZN => 
                           n11600);
   U3774 : NAND2_X1 port map( A1 => n10639, A2 => n14726, ZN => n10666);
   U3775 : XNOR2_X1 port map( A => n14450, B => n14723, ZN => n11313);
   U3776 : CLKBUF_X2 port map( A => n8330, Z => n13813);
   U3777 : AND3_X1 port map( A1 => n10746, A2 => n10837, A3 => n10836, ZN => 
                           n14927);
   U3778 : CLKBUF_X2 port map( A => n8326, Z => n10742);
   U3779 : CLKBUF_X1 port map( A => n11097, Z => n13980);
   U3780 : INV_X1 port map( A => n10724, ZN => n10725);
   U3782 : OR2_X1 port map( A1 => n11164, A2 => n14741, ZN => n14134);
   U3783 : BUF_X1 port map( A => n12639, Z => n13373);
   U3785 : CLKBUF_X1 port map( A => n8358, Z => n11312);
   U3786 : INV_X1 port map( A => n14468, ZN => n12230);
   U3787 : OR2_X1 port map( A1 => n10920, A2 => n10716, ZN => n13449);
   U3788 : OR2_X1 port map( A1 => n10716, A2 => n10682, ZN => n13448);
   U3789 : INV_X1 port map( A => n14723, ZN => n11594);
   U3790 : AND3_X1 port map( A1 => n14883, A2 => n14653, A3 => n14770, ZN => 
                           n13367);
   U3791 : CLKBUF_X2 port map( A => n8331, Z => n14117);
   U3792 : CLKBUF_X2 port map( A => n8349, Z => n13823);
   U3794 : BUF_X1 port map( A => n10871, Z => n10693);
   U3795 : CLKBUF_X1 port map( A => n11283, Z => n11971);
   U3796 : NAND2_X1 port map( A1 => n8353, A2 => n10983, ZN => n10713);
   U3797 : XNOR2_X1 port map( A => n10934, B => n10935, ZN => n13279);
   U3798 : XNOR2_X1 port map( A => n11680, B => n10647, ZN => n11570);
   U3799 : XNOR2_X1 port map( A => n11549, B => n11548, ZN => n11680);
   U3800 : NAND2_X1 port map( A1 => n11641, A2 => n11642, ZN => n11645);
   U3801 : MUX2_X2 port map( A => n13346, B => n12805, S => n10635, Z => n11366
                           );
   U3802 : XNOR2_X1 port map( A => n10648, B => n10646, ZN => n10947);
   U3803 : NAND2_X1 port map( A1 => n10708, A2 => n12992, ZN => n10648);
   U3805 : NAND2_X1 port map( A1 => intadd_46_A_3_port, A2 => 
                           intadd_46_B_3_port, ZN => n10649);
   U3806 : OAI21_X1 port map( B1 => intadd_46_B_3_port, B2 => 
                           intadd_46_A_3_port, A => intadd_46_n3, ZN => n10650)
                           ;
   U3807 : XNOR2_X1 port map( A => intadd_46_A_3_port, B => intadd_46_B_3_port,
                           ZN => n10651);
   U3808 : XNOR2_X1 port map( A => n11226, B => n10950, ZN => n11029);
   U3809 : XNOR2_X1 port map( A => n11260, B => n10652, ZN => n10896);
   U3810 : OAI211_X1 port map( C1 => n13618, C2 => n13602, A => n13616, B => 
                           n10653, ZN => n13527);
   U3811 : OAI22_X1 port map( A1 => n13618, A2 => n10653, B1 => n13620, B2 => 
                           n13619, ZN => n14748);
   U3812 : AOI21_X1 port map( B1 => n13618, B2 => n10653, A => n13616, ZN => 
                           n14752);
   U3814 : NAND2_X1 port map( A1 => n13265, A2 => n10861, ZN => n13266);
   U3815 : XNOR2_X1 port map( A => n8333, B => n10861, ZN => n11161);
   U3816 : NAND2_X1 port map( A1 => n12158, A2 => n10861, ZN => n12160);
   U3817 : XNOR2_X1 port map( A => n10656, B => n10655, ZN => n11790);
   U3818 : XNOR2_X1 port map( A => n11786, B => n11785, ZN => n10656);
   U3819 : NAND2_X1 port map( A1 => n11770, A2 => n11771, ZN => n11786);
   U3820 : INV_X1 port map( A => n11790, ZN => n11819);
   U3821 : NAND3_X1 port map( A1 => n14719, A2 => n14781, A3 => n14507, ZN => 
                           n13965);
   U3822 : INV_X1 port map( A => n12808, ZN => n10658);
   U3824 : AOI21_X2 port map( B1 => n11689, B2 => n11688, A => n11687, ZN => 
                           n14065);
   U3825 : NAND2_X1 port map( A1 => n11072, A2 => n11071, ZN => n10662);
   U3826 : NOR2_X1 port map( A1 => n10663, A2 => n12996, ZN => n12183);
   U3827 : INV_X1 port map( A => n12997, ZN => n10663);
   U3828 : NAND3_X1 port map( A1 => n12179, A2 => n12180, A3 => n12181, ZN => 
                           n10664);
   U3829 : XNOR2_X1 port map( A => n10670, B => n13408, ZN => n13410);
   U3830 : NAND2_X1 port map( A1 => n13388, A2 => n10670, ZN => n10667);
   U3831 : XNOR2_X1 port map( A => n13668, B => n13669, ZN => n10672);
   U3832 : XNOR2_X1 port map( A => n13416, B => n13417, ZN => n10673);
   U3833 : AND2_X1 port map( A1 => n14184, A2 => n14796, ZN => n10676);
   U3834 : NAND2_X1 port map( A1 => n11207, A2 => n11206, ZN => n10677);
   U3835 : BUF_X1 port map( A => intadd_66_SUM_1_port, Z => n10678);
   U3836 : INV_X1 port map( A => n14499, ZN => n10679);
   U3837 : NAND2_X1 port map( A1 => n10857, A2 => n10861, ZN => n11957);
   U3838 : XNOR2_X1 port map( A => n14441, B => EXP_out_round_7_port, ZN => 
                           n10681);
   U3839 : XNOR2_X1 port map( A => n14441, B => EXP_out_round_7_port, ZN => 
                           n12475);
   U3840 : NAND2_X1 port map( A1 => n13668, A2 => n13670, ZN => n10683);
   U3841 : NAND2_X1 port map( A1 => n13668, A2 => n13669, ZN => n10684);
   U3842 : NAND2_X1 port map( A1 => n13670, A2 => n13669, ZN => n10685);
   U3843 : NAND3_X1 port map( A1 => n10683, A2 => n10684, A3 => n10685, ZN => 
                           n13721);
   U3844 : NAND2_X1 port map( A1 => n13166, A2 => n13165, ZN => n10686);
   U3845 : INV_X1 port map( A => n14063, ZN => n10687);
   U3846 : XNOR2_X1 port map( A => n10920, B => n14478, ZN => n12135);
   U3847 : AOI22_X1 port map( A1 => n11233, A2 => n11232, B1 => n11231, B2 => 
                           n11230, ZN => n10688);
   U3848 : INV_X2 port map( A => n14465, ZN => n13914);
   U3849 : XNOR2_X1 port map( A => n10689, B => n10690, ZN => n10697);
   U3850 : XNOR2_X1 port map( A => n11657, B => n13435, ZN => n10944);
   U3851 : OAI21_X1 port map( B1 => n14121, B2 => n13236, A => n13235, ZN => 
                           n10691);
   U3852 : OR2_X1 port map( A1 => n13243, A2 => n13242, ZN => n10692);
   U3853 : BUF_X1 port map( A => n13030, Z => n10694);
   U3854 : OAI21_X1 port map( B1 => n13187, B2 => n13189, A => n13188, ZN => 
                           n10695);
   U3855 : NAND2_X1 port map( A1 => n12440, A2 => n10696, ZN => n12447);
   U3856 : INV_X1 port map( A => n10710, ZN => n13303);
   U3857 : AND2_X1 port map( A1 => n10910, A2 => n10911, ZN => n10698);
   U3858 : AOI22_X2 port map( A1 => n13034, A2 => n13033, B1 => n13032, B2 => 
                           n13031, ZN => n13558);
   U3859 : AOI21_X1 port map( B1 => n12384, B2 => n12383, A => n12382, ZN => 
                           n10699);
   U3860 : AND3_X1 port map( A1 => n13688, A2 => n13686, A3 => n13682, ZN => 
                           n10700);
   U3861 : AND3_X1 port map( A1 => n13688, A2 => n13686, A3 => n13682, ZN => 
                           n13744);
   U3862 : BUF_X1 port map( A => n12958, Z => n10701);
   U3863 : INV_X1 port map( A => n14653, ZN => n10702);
   U3864 : AND2_X1 port map( A1 => n11659, A2 => n11658, ZN => n10703);
   U3865 : OR2_X1 port map( A1 => n10704, A2 => n10864, ZN => n11119);
   U3866 : OR2_X1 port map( A1 => n13312, A2 => n13311, ZN => n10705);
   U3868 : NAND2_X1 port map( A1 => n12482, A2 => n12362, ZN => n10707);
   U3869 : XOR2_X1 port map( A => n10722, B => n10920, Z => n11371);
   U3870 : NAND2_X1 port map( A1 => n12187, A2 => n12186, ZN => n10708);
   U3871 : XNOR2_X1 port map( A => n10709, B => n11268, ZN => n10888);
   U3872 : AND2_X1 port map( A1 => n11267, A2 => n11266, ZN => n10709);
   U3873 : XNOR2_X1 port map( A => n13300, B => n10711, ZN => n10710);
   U3874 : XOR2_X1 port map( A => n13299, B => n13298, Z => n10711);
   U3876 : OR2_X2 port map( A1 => n10714, A2 => n10866, ZN => n12783);
   U3877 : XOR2_X1 port map( A => n12879, B => n12878, Z => n10715);
   U3878 : NAND2_X1 port map( A1 => n13286, A2 => n13285, ZN => n10719);
   U3879 : NAND2_X1 port map( A1 => n13286, A2 => n13285, ZN => n10720);
   U3880 : BUF_X2 port map( A => n10737, Z => n10738);
   U3881 : AND2_X1 port map( A1 => n13047, A2 => n13046, ZN => n10721);
   U3882 : XNOR2_X1 port map( A => n13277, B => n10722, ZN => n11857);
   U3883 : NAND2_X1 port map( A1 => n11563, A2 => n11562, ZN => n10723);
   U3886 : NAND2_X1 port map( A1 => n10695, A2 => n12040, ZN => n10727);
   U3887 : NAND2_X1 port map( A1 => n10707, A2 => n12563, ZN => n10728);
   U3889 : NAND2_X1 port map( A1 => n11864, A2 => n11863, ZN => n10730);
   U3890 : AOI21_X1 port map( B1 => n10681, B2 => EXP_neg, A => n12349, ZN => 
                           n10937);
   U3891 : OR2_X1 port map( A1 => n13634, A2 => n13438, ZN => n10731);
   U3892 : NAND2_X1 port map( A1 => n10731, A2 => n13437, ZN => n13440);
   U3894 : OR2_X1 port map( A1 => n10733, A2 => n14469, ZN => n11704);
   U3895 : BUF_X1 port map( A => n13312, Z => n10734);
   U3897 : XNOR2_X1 port map( A => n13091, B => n10739, ZN => n13158);
   U3898 : XNOR2_X1 port map( A => n13089, B => n13088, ZN => n10739);
   U3899 : AND2_X1 port map( A1 => n11456, A2 => n11455, ZN => n10741);
   U3900 : BUF_X1 port map( A => n12043, Z => n10744);
   U3901 : CLKBUF_X1 port map( A => n12528, Z => n14373);
   U3902 : OR2_X1 port map( A1 => n10929, A2 => n10806, ZN => n10928);
   U3904 : XNOR2_X1 port map( A => n10811, B => n10808, ZN => n14462);
   U3905 : NOR2_X1 port map( A1 => n10811, A2 => n14679, ZN => n10809);
   U3909 : OR2_X1 port map( A1 => n10818, A2 => n14553, ZN => n13708);
   U3910 : OR2_X1 port map( A1 => n10819, A2 => n12531, ZN => n13690);
   U3911 : AND2_X1 port map( A1 => n14931, A2 => n14437, ZN => n10825);
   U3912 : INV_X1 port map( A => n14768, ZN => n14518);
   U3913 : INV_X1 port map( A => I1_I1_N13, ZN => n14646);
   U3914 : INV_X1 port map( A => n14831, ZN => n14522);
   U3917 : NOR2_X1 port map( A1 => n14669, A2 => n14671, ZN => n10850);
   U3918 : NAND2_X1 port map( A1 => n14703, A2 => FP_A(21), ZN => n10851);
   U3919 : FA_X1 port map( A => n14648, B => n14649, CI => intadd_47_SUM_3_port
                           , CO => n_1338, S => n10853);
   U3920 : INV_X1 port map( A => n14662, ZN => n14454);
   U3922 : NOR2_X1 port map( A1 => FP_A(17), A2 => n14669, ZN => n10880);
   U3923 : NAND3_X2 port map( A1 => n14883, A2 => n14653, A3 => n14770, ZN => 
                           n10885);
   U3924 : NAND3_X1 port map( A1 => n14883, A2 => n14653, A3 => n14770, ZN => 
                           n10886);
   U3925 : NAND2_X1 port map( A1 => n11737, A2 => n11736, ZN => n11742);
   U3926 : AOI22_X1 port map( A1 => n13513, A2 => n13514, B1 => n13512, B2 => 
                           n13511, ZN => n13640);
   U3927 : INV_X1 port map( A => n13206, ZN => n10893);
   U3928 : INV_X1 port map( A => n11526, ZN => n11527);
   U3929 : NAND2_X1 port map( A1 => n11442, A2 => n10953, ZN => n11156);
   U3930 : INV_X1 port map( A => n11462, ZN => n10953);
   U3931 : OR2_X1 port map( A1 => n11185, A2 => n11186, ZN => n11788);
   U3932 : NAND2_X1 port map( A1 => n11185, A2 => n11186, ZN => n11787);
   U3933 : NAND2_X1 port map( A1 => n11450, A2 => n11451, ZN => n11719);
   U3934 : AOI22_X1 port map( A1 => n12902, A2 => n12901, B1 => n12938, B2 => 
                           n12900, ZN => n12909);
   U3935 : NOR2_X1 port map( A1 => FP_A(11), A2 => n14667, ZN => n10862);
   U3936 : INV_X1 port map( A => n12149, ZN => n13040);
   U3937 : NAND2_X1 port map( A1 => n13162, A2 => n10890, ZN => n11688);
   U3938 : INV_X1 port map( A => n11686, ZN => n10890);
   U3939 : XNOR2_X1 port map( A => n13065, B => n13566, ZN => n14207);
   U3941 : NAND2_X1 port map( A1 => n11569, A2 => n12962, ZN => n11678);
   U3942 : XNOR2_X1 port map( A => n13162, B => n11686, ZN => n11534);
   U3943 : INV_X1 port map( A => n13294, ZN => n10958);
   U3945 : OR2_X1 port map( A1 => n11200, A2 => n11199, ZN => n11332);
   U3946 : INV_X1 port map( A => n11511, ZN => n10897);
   U3947 : NAND2_X1 port map( A1 => n12013, A2 => n12012, ZN => n13013);
   U3948 : INV_X1 port map( A => n11785, ZN => n11171);
   U3949 : NAND2_X1 port map( A1 => n11147, A2 => n11148, ZN => n11462);
   U3950 : OR2_X1 port map( A1 => n13041, A2 => n13042, ZN => n12171);
   U3951 : AND2_X1 port map( A1 => n11612, A2 => n13058, ZN => n10965);
   U3952 : INV_X1 port map( A => n11742, ZN => n11760);
   U3953 : NAND2_X1 port map( A1 => n11417, A2 => n11416, ZN => n11526);
   U3954 : NAND2_X1 port map( A1 => n11420, A2 => n11419, ZN => n11524);
   U3955 : NOR2_X1 port map( A1 => n11423, A2 => n10972, ZN => n11528);
   U3956 : INV_X1 port map( A => n11421, ZN => n11423);
   U3957 : OR2_X1 port map( A1 => n11385, A2 => n14464, ZN => n11080);
   U3958 : INV_X1 port map( A => n13006, ZN => n13007);
   U3959 : NAND2_X1 port map( A1 => n11787, A2 => n11788, ZN => n10966);
   U3960 : OR2_X1 port map( A1 => n11188, A2 => n11187, ZN => n11811);
   U3961 : OAI21_X1 port map( B1 => n11789, B2 => n10967, A => n11788, ZN => 
                           n11813);
   U3962 : INV_X1 port map( A => n11787, ZN => n10967);
   U3963 : INV_X1 port map( A => n11691, ZN => n11474);
   U3964 : INV_X1 port map( A => n11719, ZN => n11718);
   U3965 : NOR2_X1 port map( A1 => n14435, A2 => n14509, ZN => n14436);
   U3966 : AND2_X1 port map( A1 => n11366, A2 => n11362, ZN => n10956);
   U3967 : AND2_X1 port map( A1 => n11728, A2 => n10960, ZN => n13181);
   U3970 : OR2_X1 port map( A1 => n11212, A2 => n11211, ZN => n11355);
   U3971 : NAND2_X1 port map( A1 => n10891, A2 => n11688, ZN => n13163);
   U3972 : NAND2_X1 port map( A1 => n13161, A2 => n10892, ZN => n10891);
   U3973 : NAND2_X1 port map( A1 => n10894, A2 => n11686, ZN => n10892);
   U3974 : NAND2_X1 port map( A1 => n13662, A2 => n13661, ZN => n14214);
   U3975 : NAND2_X1 port map( A1 => n13660, A2 => n13659, ZN => n13662);
   U3976 : NAND2_X1 port map( A1 => n13124, A2 => n10899, ZN => n13125);
   U3979 : NAND2_X1 port map( A1 => n11576, A2 => n13623, ZN => n11577);
   U3980 : OR2_X1 port map( A1 => n14355, A2 => n14354, ZN => n14525);
   U3981 : INV_X2 port map( A => n14653, ZN => n13809);
   U3982 : NOR2_X2 port map( A1 => n14483, A2 => n10866, ZN => n11743);
   U3983 : OR2_X1 port map( A1 => n13089, A2 => n13088, ZN => n10887);
   U3984 : INV_X1 port map( A => n13162, ZN => n10894);
   U3986 : OR2_X1 port map( A1 => n11472, A2 => n11473, ZN => n11692);
   U3987 : XNOR2_X1 port map( A => n10896, B => n11269, ZN => n10895);
   U3988 : NAND2_X1 port map( A1 => n10896, A2 => n11269, ZN => n13563);
   U3989 : XNOR2_X1 port map( A => n10888, B => n10895, ZN => n10921);
   U3990 : OR2_X1 port map( A1 => n10896, A2 => n11269, ZN => n13562);
   U3991 : NAND2_X1 port map( A1 => n10897, A2 => n11093, ZN => n11095);
   U3992 : AND2_X2 port map( A1 => n11088, A2 => n11087, ZN => n11511);
   U3993 : XNOR2_X1 port map( A => n10898, B => n13054, ZN => n13056);
   U3994 : NAND2_X1 port map( A1 => n10898, A2 => n11608, ZN => n11612);
   U3995 : OR2_X1 port map( A1 => n11608, A2 => n10898, ZN => n11613);
   U3996 : NAND2_X1 port map( A1 => n13121, A2 => n10900, ZN => n12932);
   U3997 : INV_X1 port map( A => n12913, ZN => n10899);
   U3998 : NAND2_X1 port map( A1 => n10900, A2 => n13123, ZN => n12913);
   U3999 : NAND3_X1 port map( A1 => n12908, A2 => n12909, A3 => n12907, ZN => 
                           n10900);
   U4000 : XNOR2_X1 port map( A => n13640, B => n10902, ZN => n10901);
   U4001 : INV_X1 port map( A => n13639, ZN => n10902);
   U4002 : OR2_X1 port map( A1 => n13506, A2 => n13505, ZN => n10903);
   U4003 : INV_X1 port map( A => n10921, ZN => n13579);
   U4004 : BUF_X2 port map( A => n8333, Z => n10904);
   U4006 : NAND2_X1 port map( A1 => n12155, A2 => n12153, ZN => n10907);
   U4007 : NAND2_X1 port map( A1 => n12155, A2 => n12154, ZN => n10908);
   U4008 : NAND2_X1 port map( A1 => n12153, A2 => n12154, ZN => n10909);
   U4009 : NAND3_X1 port map( A1 => n10907, A2 => n10908, A3 => n10909, ZN => 
                           n12993);
   U4010 : XNOR2_X1 port map( A => n13051, B => n11634, ZN => n12153);
   U4011 : NAND2_X1 port map( A1 => n14002, A2 => n12134, ZN => n10910);
   U4012 : NAND2_X1 port map( A1 => n12133, A2 => n12132, ZN => n10911);
   U4013 : AND2_X1 port map( A1 => n10910, A2 => n10911, ZN => n13035);
   U4014 : NAND2_X1 port map( A1 => n12781, A2 => n12782, ZN => n13295);
   U4015 : BUF_X2 port map( A => n4381, Z => n10913);
   U4016 : BUF_X2 port map( A => n4381, Z => n10914);
   U4017 : NAND2_X1 port map( A1 => n11962, A2 => n11961, ZN => n10915);
   U4018 : INV_X1 port map( A => n12925, ZN => n10916);
   U4019 : OR2_X1 port map( A1 => n14192, A2 => n14191, ZN => n10917);
   U4020 : XNOR2_X1 port map( A => n13149, B => n13148, ZN => n10918);
   U4021 : OR2_X1 port map( A1 => n13189, A2 => n13188, ZN => n10919);
   U4022 : XNOR2_X1 port map( A => n11649, B => n10920, ZN => n11222);
   U4023 : OR2_X2 port map( A1 => n10922, A2 => n10882, ZN => n13968);
   U4024 : AND2_X1 port map( A1 => n13586, A2 => n10923, ZN => n11674);
   U4025 : NAND2_X1 port map( A1 => n13585, A2 => n13587, ZN => n10923);
   U4026 : NAND2_X1 port map( A1 => n14759, A2 => n10871, ZN => n10925);
   U4027 : XOR2_X1 port map( A => n14358, B => n14357, Z => n10926);
   U4028 : NAND2_X1 port map( A1 => n12447, A2 => n12446, ZN => n10927);
   U4029 : NAND2_X1 port map( A1 => n12447, A2 => n12446, ZN => n14323);
   U4030 : OR2_X1 port map( A1 => n10929, A2 => n10806, ZN => n12488);
   U4031 : NOR2_X1 port map( A1 => n12252, A2 => n14896, ZN => n10930);
   U4032 : AND2_X1 port map( A1 => n10930, A2 => n10931, ZN => n12250);
   U4033 : AND2_X1 port map( A1 => n10932, A2 => n10942, ZN => n10931);
   U4034 : INV_X1 port map( A => n11299, ZN => n10932);
   U4036 : AOI21_X1 port map( B1 => n10681, B2 => EXP_neg, A => n12349, ZN => 
                           n10936);
   U4037 : AOI21_X1 port map( B1 => n12475, B2 => EXP_neg, A => n12349, ZN => 
                           n14931);
   U4038 : INV_X1 port map( A => n10634, ZN => n10938);
   U4039 : BUF_X2 port map( A => n14021, Z => n10939);
   U4041 : NAND2_X1 port map( A1 => n8358, A2 => n14586, ZN => n14021);
   U4043 : MUX2_X1 port map( A => n10943, B => n14471, S => n14729, Z => n10942
                           );
   U4044 : XOR2_X1 port map( A => n11672, B => n13522, Z => n10945);
   U4046 : OR2_X1 port map( A1 => n13312, A2 => n13311, ZN => n13398);
   U4047 : XOR2_X1 port map( A => n14712, B => n10948, Z => n11120);
   U4048 : NOR2_X1 port map( A1 => n11427, A2 => n11426, ZN => n10949);
   U4049 : MUX2_X1 port map( A => n11650, B => n11343, S => n10950, Z => n11345
                           );
   U4050 : MUX2_X1 port map( A => n13283, B => n14716, S => n10635, Z => n11344
                           );
   U4051 : XNOR2_X1 port map( A => n11803, B => n10951, ZN => n11804);
   U4052 : XNOR2_X1 port map( A => n11476, B => n11475, ZN => n10951);
   U4053 : NAND2_X1 port map( A1 => n13824, A2 => n10952, ZN => n12102);
   U4054 : MUX2_X1 port map( A => n13822, B => n10952, S => n14594, Z => n12633
                           );
   U4055 : MUX2_X1 port map( A => n13822, B => n10952, S => n14025, Z => n11025
                           );
   U4056 : MUX2_X1 port map( A => n13822, B => n10952, S => n10831, Z => n12710
                           );
   U4057 : MUX2_X1 port map( A => n10952, B => n13822, S => n10913, Z => n13275
                           );
   U4058 : MUX2_X1 port map( A => n10952, B => n13822, S => n8334, Z => n13826)
                           ;
   U4059 : MUX2_X1 port map( A => n10952, B => n13822, S => n10631, Z => n12651
                           );
   U4060 : MUX2_X1 port map( A => n10952, B => n13822, S => n13450, Z => n12239
                           );
   U4061 : MUX2_X1 port map( A => n10952, B => n13822, S => n8351, Z => n11656)
                           ;
   U4062 : MUX2_X1 port map( A => n13822, B => n10952, S => n14945, Z => n12786
                           );
   U4063 : MUX2_X1 port map( A => n10952, B => n13822, S => n11738, Z => n11285
                           );
   U4064 : MUX2_X1 port map( A => n10952, B => n13822, S => n10635, Z => n11872
                           );
   U4065 : MUX2_X1 port map( A => n10952, B => n13822, S => n13364, Z => n12737
                           );
   U4066 : MUX2_X1 port map( A => n10952, B => n13822, S => n13327, Z => n13330
                           );
   U4067 : MUX2_X1 port map( A => n10952, B => n13822, S => n13261, Z => n12199
                           );
   U4068 : MUX2_X1 port map( A => n10952, B => n13822, S => n10742, Z => n13246
                           );
   U4069 : MUX2_X1 port map( A => n10952, B => n13822, S => n11703, Z => n11255
                           );
   U4070 : MUX2_X1 port map( A => n10952, B => n13822, S => n13813, Z => n12722
                           );
   U4071 : MUX2_X1 port map( A => n13822, B => n10952, S => n10841, Z => n12215
                           );
   U4072 : MUX2_X1 port map( A => n10952, B => n13822, S => n8329, Z => n12662)
                           ;
   U4073 : NAND2_X1 port map( A1 => n12163, A2 => n10952, ZN => n12631);
   U4074 : NAND2_X1 port map( A1 => n11476, A2 => n11475, ZN => n11800);
   U4075 : OR2_X1 port map( A1 => n11476, A2 => n11475, ZN => n11801);
   U4076 : NAND2_X1 port map( A1 => n13091, A2 => n13090, ZN => n10954);
   U4077 : NAND2_X1 port map( A1 => n10887, A2 => n10954, ZN => n13104);
   U4078 : NAND3_X1 port map( A1 => n10954, A2 => n10887, A3 => n13102, ZN => 
                           n13152);
   U4079 : NAND2_X1 port map( A1 => n11366, A2 => n10955, ZN => n11368);
   U4080 : XNOR2_X1 port map( A => n13883, B => n10956, ZN => intadd_66_CI);
   U4081 : INV_X1 port map( A => n13295, ZN => n12788);
   U4082 : OR2_X1 port map( A1 => n11126, A2 => n11142, ZN => n11215);
   U4083 : AOI22_X1 port map( A1 => n10959, A2 => n14363, B1 => n14361, B2 => 
                           n14362, ZN => n14907);
   U4084 : NAND2_X1 port map( A1 => n10926, A2 => n14359, ZN => n10959);
   U4085 : NAND2_X1 port map( A1 => n13180, A2 => n13181, ZN => n11735);
   U4088 : XNOR2_X1 port map( A => n10976, B => n14775, ZN => n14762);
   U4089 : NAND2_X1 port map( A1 => n10964, A2 => n10963, ZN => n14775);
   U4090 : NAND2_X1 port map( A1 => n11683, A2 => n11682, ZN => n10963);
   U4091 : OAI21_X1 port map( B1 => n11683, B2 => n11682, A => n11681, ZN => 
                           n10964);
   U4092 : NAND3_X1 port map( A1 => n11610, A2 => n11609, A3 => n10965, ZN => 
                           n13569);
   U4093 : NAND2_X1 port map( A1 => n14210, A2 => n10889, ZN => n14830);
   U4096 : OR2_X1 port map( A1 => n14257, A2 => n13658, ZN => n13661);
   U4097 : NAND2_X1 port map( A1 => n14257, A2 => n13658, ZN => n13659);
   U4098 : OR2_X1 port map( A1 => n13292, A2 => n13291, ZN => n13313);
   U4099 : AND3_X1 port map( A1 => n14605, A2 => FP_A(7), A3 => FP_A(8), ZN => 
                           n10865);
   U4100 : AND2_X1 port map( A1 => n12634, A2 => n12633, ZN => n13091);
   U4101 : XNOR2_X1 port map( A => n12924, B => n12923, ZN => n13128);
   U4102 : OR2_X1 port map( A1 => n11336, A2 => n10677, ZN => n11337);
   U4104 : AOI22_X1 port map( A1 => n11499, A2 => n11498, B1 => n11497, B2 => 
                           n11496, ZN => n11507);
   U4105 : XNOR2_X1 port map( A => n13135, B => n13134, ZN => n13216);
   U4106 : OR2_X1 port map( A1 => n11020, A2 => n11019, ZN => n11072);
   U4107 : OAI22_X1 port map( A1 => n13723, A2 => n13722, B1 => n13721, B2 => 
                           n13720, ZN => n13728);
   U4109 : XNOR2_X1 port map( A => n11919, B => n14085, ZN => n13221);
   U4110 : NOR2_X1 port map( A1 => n11830, A2 => n11829, ZN => n11832);
   U4111 : XNOR2_X1 port map( A => n13133, B => n13132, ZN => n13135);
   U4112 : NAND2_X1 port map( A1 => n12043, A2 => n12042, ZN => n12044);
   U4113 : OAI211_X1 port map( C1 => n10916, C2 => n13127, A => n13126, B => 
                           n13125, ZN => n13215);
   U4114 : OR2_X1 port map( A1 => n11636, A2 => n11635, ZN => n12151);
   U4115 : OR2_X1 port map( A1 => n11427, A2 => n11426, ZN => n11544);
   U4117 : XNOR2_X1 port map( A => n11575, B => n11683, ZN => n13626);
   U4118 : INV_X1 port map( A => n11676, ZN => n11677);
   U4119 : OR2_X1 port map( A1 => n11243, A2 => n11241, ZN => n11670);
   U4120 : XNOR2_X1 port map( A => n14084, B => n14083, ZN => n11919);
   U4121 : NAND2_X1 port map( A1 => n14783, A2 => n10871, ZN => n14118);
   U4122 : OR2_X1 port map( A1 => n13868, A2 => n10913, ZN => n10968);
   U4123 : OR2_X1 port map( A1 => n13868, A2 => n10973, ZN => n10969);
   U4124 : INV_X1 port map( A => n14256, ZN => n13658);
   U4125 : NAND2_X1 port map( A1 => n12101, A2 => n12342, ZN => n10970);
   U4127 : AND2_X1 port map( A1 => n14460, A2 => n14783, ZN => n10971);
   U4128 : AND2_X1 port map( A1 => n11422, A2 => n14727, ZN => n10972);
   U4129 : AND2_X1 port map( A1 => n11167, A2 => n11166, ZN => n10974);
   U4131 : XNOR2_X1 port map( A => n11359, B => n12260, ZN => n12043);
   U4132 : XOR2_X1 port map( A => n12233, B => n14065, Z => n10976);
   U4133 : AND2_X1 port map( A1 => n12124, A2 => n14488, ZN => n10977);
   U4134 : INV_X1 port map( A => n13885, ZN => n11406);
   U4135 : NAND2_X1 port map( A1 => n11473, A2 => n11472, ZN => n11691);
   U4136 : NAND2_X1 port map( A1 => n13967, A2 => n14735, ZN => n11248);
   U4137 : NOR2_X1 port map( A1 => n11305, A2 => n14841, ZN => n11492);
   U4138 : INV_X1 port map( A => n13013, ZN => n13014);
   U4139 : NAND2_X1 port map( A1 => n11170, A2 => n11169, ZN => n11785);
   U4140 : NAND2_X1 port map( A1 => n14725, A2 => n10864, ZN => n11707);
   U4141 : XNOR2_X1 port map( A => n11552, B => n11551, ZN => n11554);
   U4142 : NAND2_X1 port map( A1 => n12027, A2 => n13002, ZN => n13006);
   U4143 : OR2_X1 port map( A1 => n11786, A2 => n10974, ZN => n11172);
   U4144 : INV_X1 port map( A => n11248, ZN => n14002);
   U4145 : OAI21_X1 port map( B1 => n11717, B2 => n12866, A => n12864, ZN => 
                           n11792);
   U4146 : NAND2_X1 port map( A1 => n11652, A2 => n11649, ZN => n11653);
   U4147 : XNOR2_X1 port map( A => n11554, B => n11553, ZN => n11565);
   U4148 : NAND2_X1 port map( A1 => n11850, A2 => n11849, ZN => n13028);
   U4149 : MUX2_X1 port map( A => n11385, B => n11933, S => n10869, Z => n11937
                           );
   U4150 : XNOR2_X1 port map( A => n13426, B => n13629, ZN => n11664);
   U4151 : INV_X1 port map( A => n13028, ZN => n12995);
   U4152 : AND2_X1 port map( A1 => n13042, A2 => n13041, ZN => n12172);
   U4153 : BUF_X1 port map( A => n8330, Z => n13810);
   U4154 : OAI211_X1 port map( C1 => n13346, C2 => n8329, A => n11654, B => 
                           n11653, ZN => n13433);
   U4155 : XNOR2_X1 port map( A => n12922, B => n12921, ZN => n12924);
   U4157 : XNOR2_X1 port map( A => n11664, B => n13630, ZN => n11666);
   U4158 : BUF_X1 port map( A => n14653, Z => n13482);
   U4160 : OR2_X1 port map( A1 => n13727, A2 => n13302, ZN => n13305);
   U4161 : XNOR2_X1 port map( A => n12035, B => n12034, ZN => n13144);
   U4162 : XNOR2_X1 port map( A => n11543, B => n11542, ZN => n12957);
   U4163 : XNOR2_X1 port map( A => n12624, B => n12623, ZN => n13156);
   U4164 : NAND2_X1 port map( A1 => n11679, A2 => n11548, ZN => n11108);
   U4165 : NAND2_X1 port map( A1 => n13731, A2 => n13744, ZN => n12528);
   U4168 : NAND2_X1 port map( A1 => n13642, A2 => n13641, ZN => n14257);
   U4169 : NAND2_X1 port map( A1 => n11109, A2 => n11108, ZN => n11684);
   U4170 : INV_X1 port map( A => n11678, ZN => n11682);
   U4171 : OAI21_X1 port map( B1 => n12043, B2 => n12042, A => intadd_66_n2, ZN
                           => n12045);
   U4172 : NAND2_X1 port map( A1 => n11482, A2 => n11481, ZN => n14755);
   U4173 : NAND2_X1 port map( A1 => n12045, A2 => n12044, ZN => intadd_66_n1);
   U4174 : OAI21_X1 port map( B1 => n11833, B2 => n11832, A => n11831, ZN => 
                           n14801);
   U4178 : MUX2_X1 port map( A => n14833, B => n12783, S => n13327, Z => n10980
                           );
   U4179 : XOR2_X1 port map( A => n10914, B => n14725, Z => n10978);
   U4180 : NAND2_X1 port map( A1 => n10978, A2 => n14727, ZN => n10979);
   U4181 : AND2_X1 port map( A1 => n10980, A2 => n10979, ZN => n13071);
   U4182 : NAND2_X1 port map( A1 => n14778, A2 => n14720, ZN => n11418);
   U4183 : BUF_X2 port map( A => n11418, Z => n14017);
   U4184 : MUX2_X1 port map( A => n11900, B => n11201, S => n13823, Z => n10982
                           );
   U4185 : INV_X1 port map( A => n14484, ZN => n13915);
   U4186 : MUX2_X1 port map( A => n13915, B => n14779, S => n13282, Z => n10981
                           );
   U4187 : XNOR2_X1 port map( A => n13071, B => n13073, ZN => n10986);
   U4188 : MUX2_X1 port map( A => n14114, B => n13362, S => n13924, Z => n10985
                           );
   U4189 : AND2_X1 port map( A1 => n384, A2 => n14602, ZN => n10875);
   U4190 : NOR2_X1 port map( A1 => n14601, A2 => FP_A(17), ZN => n10834);
   U4191 : MUX2_X1 port map( A => n12146, B => n11225, S => n8401, Z => n10984)
                           ;
   U4192 : XNOR2_X1 port map( A => n10986, B => n13072, ZN => n10997);
   U4193 : NAND2_X2 port map( A1 => n8338, A2 => n14736, ZN => n13868);
   U4194 : MUX2_X1 port map( A => n10640, B => n13868, S => n14477, Z => n10989
                           );
   U4195 : XNOR2_X1 port map( A => n12124, B => n10869, ZN => n10987);
   U4196 : NAND2_X1 port map( A1 => n14813, A2 => n10987, ZN => n10988);
   U4197 : NAND2_X1 port map( A1 => n10989, A2 => n10988, ZN => n12894);
   U4198 : NAND3_X1 port map( A1 => FP_A(3), A2 => FP_A(4), A3 => n14596, ZN =>
                           n10881);
   U4199 : MUX2_X1 port map( A => n14728, B => n13980, S => n13813, Z => n10992
                           );
   U4200 : INV_X2 port map( A => n14721, ZN => n12014);
   U4201 : XNOR2_X1 port map( A => n8329, B => n12014, ZN => n10990);
   U4202 : NAND2_X1 port map( A1 => n14786, A2 => n10990, ZN => n10991);
   U4204 : XNOR2_X1 port map( A => n12894, B => n12895, ZN => n10995);
   U4205 : NAND2_X2 port map( A1 => n14780, A2 => n14713, ZN => n13371);
   U4206 : MUX2_X1 port map( A => n13372, B => n13371, S => B_SIG_8_port, Z => 
                           n10994);
   U4207 : NAND3_X1 port map( A1 => FP_A(15), A2 => n14580, A3 => n14661, ZN =>
                           n10883);
   U4208 : MUX2_X1 port map( A => n13373, B => n10745, S => n13485, Z => n10993
                           );
   U4210 : XNOR2_X1 port map( A => n10995, B => n12906, ZN => n10996);
   U4211 : NAND2_X1 port map( A1 => n10997, A2 => n10996, ZN => n12934);
   U4212 : NAND2_X1 port map( A1 => n12935, A2 => n12934, ZN => n11023);
   U4213 : NAND2_X1 port map( A1 => n14759, A2 => n14777, ZN => n10998);
   U4214 : NAND2_X1 port map( A1 => n10998, A2 => n10693, ZN => n11002);
   U4215 : BUF_X2 port map( A => n11321, Z => n11226);
   U4216 : NAND2_X1 port map( A1 => n14711, A2 => n14594, ZN => n10999);
   U4218 : OAI21_X1 port map( B1 => n11226, B2 => n10999, A => n13277, ZN => 
                           n11001);
   U4219 : BUF_X4 port map( A => n381, Z => n14025);
   U4220 : XNOR2_X1 port map( A => n13277, B => n14025, ZN => n11000);
   U4221 : AOI22_X1 port map( A1 => n11002, A2 => n11001, B1 => n13279, B2 => 
                           n11000, ZN => n11006);
   U4222 : NAND2_X1 port map( A1 => n14789, A2 => n14719, ZN => n11007);
   U4223 : NAND2_X1 port map( A1 => n11006, A2 => n11007, ZN => n11066);
   U4224 : NAND2_X1 port map( A1 => n14741, A2 => n14787, ZN => n11013);
   U4225 : BUF_X2 port map( A => n11013, Z => n13283);
   U4226 : MUX2_X1 port map( A => n13283, B => n14716, S => n13485, Z => n11005
                           );
   U4227 : XNOR2_X1 port map( A => n8340, B => n14584, ZN => n11237);
   U4228 : XNOR2_X1 port map( A => n11703, B => n10877, ZN => n11003);
   U4229 : NAND2_X1 port map( A1 => n11005, A2 => n11004, ZN => n11067);
   U4230 : NAND2_X1 port map( A1 => n11066, A2 => n11067, ZN => n11010);
   U4231 : INV_X1 port map( A => n11006, ZN => n11009);
   U4232 : INV_X1 port map( A => n11007, ZN => n11008);
   U4233 : NAND2_X1 port map( A1 => n11009, A2 => n11008, ZN => n11065);
   U4234 : NAND2_X1 port map( A1 => n11010, A2 => n11065, ZN => n11073);
   U4235 : NAND2_X1 port map( A1 => n14454, A2 => FP_A(7), ZN => n10856);
   U4236 : MUX2_X1 port map( A => n11043, B => n10680, S => n13234, Z => n11012
                           );
   U4237 : NAND2_X1 port map( A1 => n14724, A2 => n14710, ZN => n10860);
   U4238 : BUF_X2 port map( A => n11149, Z => n11834);
   U4239 : MUX2_X1 port map( A => n10725, B => n11149, S => n14449, Z => n11011
                           );
   U4240 : NAND2_X1 port map( A1 => n11012, A2 => n11011, ZN => n13093);
   U4241 : MUX2_X1 port map( A => n13347, B => n14716, S => B_SIG_8_port, Z => 
                           n11016);
   U4242 : XNOR2_X1 port map( A => n12764, B => n11861, ZN => n11014);
   U4243 : NAND2_X1 port map( A1 => n11014, A2 => n12174, ZN => n11015);
   U4244 : NAND2_X1 port map( A1 => n11016, A2 => n11015, ZN => n13092);
   U4245 : XNOR2_X1 port map( A => n13092, B => n13093, ZN => n11020);
   U4246 : INV_X1 port map( A => n10866, ZN => n13265);
   U4247 : MUX2_X1 port map( A => n11743, B => n13323, S => n10742, Z => n11018
                           );
   U4248 : OAI21_X1 port map( B1 => n10640, B2 => n14455, A => n10968, ZN => 
                           n11017);
   U4249 : NOR2_X1 port map( A1 => n11018, A2 => n11017, ZN => n11019);
   U4250 : NAND2_X1 port map( A1 => n11020, A2 => n11019, ZN => n11071);
   U4251 : NAND2_X1 port map( A1 => n11073, A2 => n11071, ZN => n11021);
   U4252 : NAND2_X1 port map( A1 => n11021, A2 => n11072, ZN => n12933);
   U4253 : INV_X1 port map( A => n12933, ZN => n11022);
   U4254 : XNOR2_X1 port map( A => n11023, B => n11022, ZN => n11830);
   U4256 : NAND2_X2 port map( A1 => n14789, A2 => n14715, ZN => n13822);
   U4257 : BUF_X1 port map( A => n14878, Z => n13824);
   U4258 : NOR2_X1 port map( A1 => FP_A(20), A2 => n14673, ZN => n10878);
   U4259 : NAND2_X1 port map( A1 => n14722, A2 => n10878, ZN => n10870);
   U4260 : MUX2_X1 port map( A => n13824, B => n11971, S => n14594, Z => n11024
                           );
   U4261 : AND2_X1 port map( A1 => n11025, A2 => n11024, ZN => n12940);
   U4262 : MUX2_X1 port map( A => n13347, B => n14716, S => n12764, Z => n12898
                           );
   U4263 : INV_X1 port map( A => n14464, ZN => n11272);
   U4264 : XNOR2_X1 port map( A => n11272, B => n11861, ZN => n11026);
   U4265 : NAND2_X1 port map( A1 => n11026, A2 => n12174, ZN => n12897);
   U4266 : AND2_X1 port map( A1 => n12898, A2 => n12897, ZN => n12938);
   U4267 : XNOR2_X1 port map( A => n12940, B => n12938, ZN => n11039);
   U4268 : MUX2_X1 port map( A => n13449, B => n13448, S => n13327, Z => n11028
                           );
   U4269 : MUX2_X1 port map( A => n14833, B => n13451, S => n11272, Z => n11027
                           );
   U4270 : AND2_X1 port map( A1 => n11028, A2 => n11027, ZN => n12622);
   U4271 : NAND2_X1 port map( A1 => n11029, A2 => n14479, ZN => n11032);
   U4272 : MUX2_X1 port map( A => n12146, B => n11225, S => n10635, Z => n11030
                           );
   U4273 : INV_X1 port map( A => n11030, ZN => n11031);
   U4274 : NAND2_X1 port map( A1 => n11032, A2 => n11031, ZN => n11037);
   U4275 : MUX2_X1 port map( A => n13920, B => n14728, S => n10831, Z => n11035
                           );
   U4276 : XNOR2_X1 port map( A => n13813, B => n12014, ZN => n11033);
   U4277 : NAND2_X1 port map( A1 => n14786, A2 => n11033, ZN => n11034);
   U4278 : NAND2_X1 port map( A1 => n11035, A2 => n11034, ZN => n11036);
   U4279 : NAND2_X1 port map( A1 => n11037, A2 => n11036, ZN => n12620);
   U4280 : NAND2_X1 port map( A1 => n12622, A2 => n12620, ZN => n11038);
   U4281 : NAND2_X1 port map( A1 => n11038, A2 => n12621, ZN => n12942);
   U4282 : XNOR2_X1 port map( A => n11039, B => n12942, ZN => n11053);
   U4283 : MUX2_X1 port map( A => n10925, B => n10736, S => n14593, Z => n11042
                           );
   U4284 : INV_X1 port map( A => FP_B(4), ZN => n10835);
   U4285 : XOR2_X1 port map( A => n13277, B => n10635, Z => n11040);
   U4286 : NAND2_X1 port map( A1 => n10971, A2 => n11040, ZN => n11041);
   U4287 : AND2_X1 port map( A1 => n11042, A2 => n11041, ZN => n12901);
   U4288 : NAND3_X1 port map( A1 => n14883, A2 => n14770, A3 => n14719, ZN => 
                           n12900);
   U4289 : XNOR2_X1 port map( A => n12901, B => n12900, ZN => n12939);
   U4290 : MUX2_X1 port map( A => n10680, B => n11043, S => n10831, Z => n11045
                           );
   U4292 : MUX2_X1 port map( A => n10725, B => n11834, S => n12246, Z => n11044
                           );
   U4293 : NAND2_X1 port map( A1 => n11045, A2 => n11044, ZN => n11051);
   U4294 : INV_X1 port map( A => n11051, ZN => n11049);
   U4295 : MUX2_X1 port map( A => n14020, B => n10940, S => n13261, Z => n11047
                           );
   U4296 : NAND2_X1 port map( A1 => n14771, A2 => n14467, ZN => n11046);
   U4297 : NAND2_X1 port map( A1 => n11047, A2 => n11046, ZN => n11050);
   U4298 : INV_X1 port map( A => n11050, ZN => n11048);
   U4299 : NAND2_X1 port map( A1 => n11049, A2 => n11048, ZN => n12911);
   U4300 : NAND2_X1 port map( A1 => n11051, A2 => n11050, ZN => n12910);
   U4301 : NAND2_X1 port map( A1 => n12911, A2 => n12910, ZN => n12941);
   U4302 : XNOR2_X1 port map( A => n12939, B => n12941, ZN => n11052);
   U4303 : XNOR2_X1 port map( A => n11053, B => n11052, ZN => n11829);
   U4304 : INV_X1 port map( A => n11829, ZN => n11054);
   U4305 : XNOR2_X1 port map( A => n14946, B => n11054, ZN => n11110);
   U4306 : MUX2_X1 port map( A => n10640, B => n13868, S => n14457, Z => n11058
                           );
   U4307 : XOR2_X1 port map( A => n10914, B => n12124, Z => n11056);
   U4308 : NAND2_X1 port map( A1 => n14813, A2 => n11056, ZN => n11057);
   U4309 : NAND2_X1 port map( A1 => n11058, A2 => n11057, ZN => n13847);
   U4310 : MUX2_X1 port map( A => n14833, B => n12783, S => n12764, Z => n11061
                           );
   U4311 : XNOR2_X1 port map( A => n12018, B => n13328, ZN => n11059);
   U4312 : NAND2_X1 port map( A1 => n11059, A2 => n14727, ZN => n11060);
   U4313 : NAND2_X1 port map( A1 => n11061, A2 => n11060, ZN => n13852);
   U4314 : XNOR2_X1 port map( A => n13852, B => n13847, ZN => n11064);
   U4315 : MUX2_X1 port map( A => n14017, B => n11201, S => n11649, Z => n11063
                           );
   U4316 : MUX2_X1 port map( A => n13915, B => n14779, S => n13813, Z => n11062
                           );
   U4317 : NAND2_X1 port map( A1 => n11063, A2 => n11062, ZN => n13848);
   U4318 : XNOR2_X1 port map( A => n11064, B => n13848, ZN => n11571);
   U4319 : NAND2_X1 port map( A1 => n11066, A2 => n11065, ZN => n11068);
   U4320 : XNOR2_X1 port map( A => n11068, B => n11067, ZN => n11573);
   U4321 : NOR2_X1 port map( A1 => n11571, A2 => n11573, ZN => n11070);
   U4322 : NAND2_X1 port map( A1 => n11571, A2 => n11573, ZN => n11069);
   U4323 : OAI21_X1 port map( B1 => intadd_46_SUM_0_port, B2 => n11070, A => 
                           n11069, ZN => n11685);
   U4324 : MUX2_X1 port map( A => n14833, B => n12783, S => n11703, Z => n11076
                           );
   U4325 : XNOR2_X1 port map( A => n12018, B => n11738, ZN => n11074);
   U4326 : NAND2_X1 port map( A1 => n11074, A2 => n14727, ZN => n11075);
   U4327 : NAND2_X1 port map( A1 => n11076, A2 => n11075, ZN => n11521);
   U4328 : INV_X1 port map( A => n11521, ZN => n11084);
   U4329 : MUX2_X1 port map( A => n11043, B => n10680, S => n10743, Z => n11078
                           );
   U4330 : MUX2_X1 port map( A => n10725, B => n11834, S => n10914, Z => n11077
                           );
   U4331 : NAND2_X1 port map( A1 => n11078, A2 => n11077, ZN => n11522);
   U4332 : INV_X1 port map( A => n11522, ZN => n11083);
   U4333 : NAND2_X1 port map( A1 => n11522, A2 => n11521, ZN => n11082);
   U4334 : NAND2_X1 port map( A1 => n14760, A2 => n8338, ZN => n13228);
   U4335 : OR2_X1 port map( A1 => n13228, A2 => n14717, ZN => n12127);
   U4336 : NAND2_X1 port map( A1 => n12127, A2 => n14464, ZN => n11081);
   U4337 : BUF_X2 port map( A => n10866, Z => n12010);
   U4338 : XNOR2_X1 port map( A => n12010, B => n13273, ZN => n11079);
   U4339 : AOI22_X1 port map( A1 => n11081, A2 => n11080, B1 => n14813, B2 => 
                           n11079, ZN => n11519);
   U4340 : AOI22_X1 port map( A1 => n11084, A2 => n11083, B1 => n11082, B2 => 
                           n11519, ZN => n11679);
   U4341 : XNOR2_X1 port map( A => n11321, B => n14593, ZN => n11085);
   U4342 : NAND2_X1 port map( A1 => n11085, A2 => n14479, ZN => n11088);
   U4343 : OR2_X1 port map( A1 => n12146, A2 => n14447, ZN => n11086);
   U4344 : OAI21_X1 port map( B1 => n11225, B2 => n14025, A => n11086, ZN => 
                           n11087);
   U4345 : MUX2_X1 port map( A => n10925, B => n10736, S => n10864, Z => n11090
                           );
   U4346 : XNOR2_X1 port map( A => n13277, B => n14594, ZN => n11089);
   U4347 : NAND2_X1 port map( A1 => n13279, A2 => n11089, ZN => n11514);
   U4348 : NAND2_X1 port map( A1 => n11090, A2 => n11514, ZN => n11093);
   U4349 : NAND2_X1 port map( A1 => n12230, A2 => n14450, ZN => n11091);
   U4351 : INV_X1 port map( A => n11093, ZN => n11094);
   U4352 : AOI22_X1 port map( A1 => n11095, A2 => n11510, B1 => n11094, B2 => 
                           n11511, ZN => n11548);
   U4353 : NAND2_X1 port map( A1 => n14541, A2 => n14702, ZN => n10872);
   U4354 : NOR2_X1 port map( A1 => n11248, A2 => n11487, ZN => n11127);
   U4355 : MUX2_X1 port map( A => n11096, B => n13908, S => n12246, Z => n11100
                           );
   U4356 : MUX2_X1 port map( A => n13920, B => n14728, S => n10869, Z => n11098
                           );
   U4357 : INV_X1 port map( A => n11098, ZN => n11099);
   U4358 : MUX2_X1 port map( A => n13372, B => n13371, S => n8401, Z => n11102)
                           ;
   U4359 : MUX2_X1 port map( A => n10745, B => n13373, S => n14465, Z => n11101
                           );
   U4360 : NAND2_X1 port map( A1 => n11102, A2 => n11101, ZN => n11551);
   U4361 : NAND2_X1 port map( A1 => n11553, A2 => n11551, ZN => n11107);
   U4362 : BUF_X1 port map( A => n8330, Z => n13239);
   U4363 : MUX2_X1 port map( A => n11900, B => n11201, S => n13239, Z => n11104
                           );
   U4364 : MUX2_X1 port map( A => n14779, B => n14456, S => n10831, Z => n11103
                           );
   U4365 : AND2_X1 port map( A1 => n11104, A2 => n11103, ZN => n11550);
   U4366 : INV_X1 port map( A => n11553, ZN => n11106);
   U4367 : INV_X1 port map( A => n11551, ZN => n11105);
   U4368 : OAI21_X1 port map( B1 => n11679, B2 => n11548, A => n11549, ZN => 
                           n11109);
   U4369 : XNOR2_X1 port map( A => n11110, B => n11828, ZN => n13214);
   U4370 : MUX2_X1 port map( A => n11043, B => n10680, S => n11738, Z => n11112
                           );
   U4371 : MUX2_X1 port map( A => n10725, B => n11149, S => n11703, Z => n11111
                           );
   U4372 : NAND2_X1 port map( A1 => n11112, A2 => n11111, ZN => n11144);
   U4373 : MUX2_X1 port map( A => n13347, B => n14716, S => n14447, Z => n11115
                           );
   U4374 : XNOR2_X1 port map( A => n14463, B => n14593, ZN => n11113);
   U4375 : NAND2_X1 port map( A1 => n12174, A2 => n11113, ZN => n11114);
   U4376 : NAND2_X1 port map( A1 => n11115, A2 => n11114, ZN => n11145);
   U4377 : AND2_X1 port map( A1 => n11144, A2 => n11145, ZN => n11142);
   U4378 : MUX2_X1 port map( A => n14020, B => n10940, S => n13234, Z => n11117
                           );
   U4379 : NAND2_X1 port map( A1 => n14771, A2 => n14945, ZN => n11116);
   U4380 : AND2_X1 port map( A1 => n11117, A2 => n11116, ZN => n11175);
   U4381 : NAND2_X1 port map( A1 => n12142, A2 => n10864, ZN => n11118);
   U4382 : NAND2_X1 port map( A1 => n11119, A2 => n11118, ZN => n11122);
   U4383 : NAND2_X1 port map( A1 => n12640, A2 => n11120, ZN => n11121);
   U4384 : NAND2_X1 port map( A1 => n11122, A2 => n11121, ZN => n11174);
   U4385 : OAI21_X1 port map( B1 => n11861, B2 => n10884, A => n14712, ZN => 
                           n14129);
   U4387 : NAND2_X1 port map( A1 => n11174, A2 => n11173, ZN => n11125);
   U4388 : INV_X1 port map( A => n11174, ZN => n11124);
   U4389 : INV_X1 port map( A => n11173, ZN => n11123);
   U4390 : AOI22_X1 port map( A1 => n11175, A2 => n11125, B1 => n11124, B2 => 
                           n11123, ZN => n11126);
   U4391 : NAND2_X1 port map( A1 => n11142, A2 => n11126, ZN => n11213);
   U4392 : AND2_X1 port map( A1 => n11213, A2 => n11215, ZN => n11141);
   U4393 : MUX2_X1 port map( A => n11096, B => n12837, S => n11965, Z => n11130
                           );
   U4394 : MUX2_X1 port map( A => n14728, B => n13920, S => n8351, Z => n11128)
                           ;
   U4395 : INV_X1 port map( A => n11128, ZN => n11129);
   U4396 : MUX2_X1 port map( A => n14017, B => n13984, S => n10743, Z => n11132
                           );
   U4397 : MUX2_X1 port map( A => n13915, B => n14779, S => n10913, Z => n11131
                           );
   U4398 : NAND2_X1 port map( A1 => n11132, A2 => n11131, ZN => n11137);
   U4399 : NAND2_X1 port map( A1 => n11136, A2 => n11137, ZN => n11435);
   U4400 : MUX2_X1 port map( A => n13449, B => n13448, S => n14731, Z => n11135
                           );
   U4401 : MUX2_X1 port map( A => n14833, B => n13451, S => n10635, Z => n11134
                           );
   U4402 : AND2_X1 port map( A1 => n11135, A2 => n11134, ZN => n11437);
   U4403 : NAND2_X1 port map( A1 => n11435, A2 => n11437, ZN => n11140);
   U4404 : INV_X1 port map( A => n11136, ZN => n11139);
   U4405 : INV_X1 port map( A => n11137, ZN => n11138);
   U4406 : NAND2_X1 port map( A1 => n11139, A2 => n11138, ZN => n11436);
   U4407 : NAND2_X1 port map( A1 => n11140, A2 => n11436, ZN => n11214);
   U4408 : XNOR2_X1 port map( A => n11141, B => n11214, ZN => n11192);
   U4409 : INV_X1 port map( A => n11142, ZN => n11143);
   U4410 : OAI21_X1 port map( B1 => n11145, B2 => n11144, A => n11143, ZN => 
                           n11446);
   U4411 : MUX2_X1 port map( A => n13283, B => n14716, S => n14777, Z => n11148
                           );
   U4412 : XNOR2_X1 port map( A => n14463, B => n14025, ZN => n11146);
   U4413 : NAND2_X1 port map( A1 => n12174, A2 => n11146, ZN => n11147);
   U4414 : NAND2_X1 port map( A1 => n11149, A2 => n8333, ZN => n11151);
   U4415 : NAND2_X1 port map( A1 => n14451, A2 => n14818, ZN => n11150);
   U4416 : NAND2_X1 port map( A1 => n11151, A2 => n11150, ZN => n11155);
   U4417 : NAND2_X1 port map( A1 => n10857, A2 => n11152, ZN => n11154);
   U4418 : NAND2_X1 port map( A1 => n11155, A2 => n11154, ZN => n11461);
   U4419 : AND2_X1 port map( A1 => n12640, A2 => n14719, ZN => n11460);
   U4420 : NAND2_X1 port map( A1 => n11461, A2 => n11460, ZN => n11442);
   U4421 : INV_X1 port map( A => n11460, ZN => n11153);
   U4422 : NAND3_X1 port map( A1 => n11155, A2 => n11154, A3 => n11153, ZN => 
                           n11441);
   U4423 : NAND2_X1 port map( A1 => n11156, A2 => n11441, ZN => n11159);
   U4424 : MUX2_X1 port map( A => n11743, B => n13323, S => n10905, Z => n11158
                           );
   U4425 : OAI21_X1 port map( B1 => n10640, B2 => n14788, A => n10969, ZN => 
                           n11157);
   U4426 : NOR2_X1 port map( A1 => n11158, A2 => n11157, ZN => n11440);
   U4427 : OAI21_X1 port map( B1 => n11446, B2 => n11159, A => n11440, ZN => 
                           n11191);
   U4428 : NAND2_X1 port map( A1 => n11446, A2 => n11159, ZN => n11190);
   U4429 : AND2_X1 port map( A1 => n11191, A2 => n11190, ZN => n11160);
   U4430 : NAND2_X1 port map( A1 => n11192, A2 => n11160, ZN => n11431);
   U4431 : MUX2_X1 port map( A => n14818, B => n11149, S => n8352, Z => n11163)
                           ;
   U4432 : NAND2_X1 port map( A1 => n10857, A2 => n11161, ZN => n11162);
   U4433 : NAND2_X1 port map( A1 => n11163, A2 => n11162, ZN => n11770);
   U4434 : NAND2_X1 port map( A1 => n13347, A2 => n14719, ZN => n11165);
   U4435 : NOR2_X1 port map( A1 => FP_A(11), A2 => n14580, ZN => n10876);
   U4436 : AND2_X1 port map( A1 => n11165, A2 => n14134, ZN => n11771);
   U4437 : MUX2_X1 port map( A => n14017, B => n13984, S => n10914, Z => n11167
                           );
   U4438 : MUX2_X1 port map( A => n13915, B => n14779, S => n12743, Z => n11166
                           );
   U4439 : MUX2_X1 port map( A => n10640, B => n13868, S => n14448, Z => n11170
                           );
   U4440 : XOR2_X1 port map( A => n8352, B => n13265, Z => n11168);
   U4441 : NAND2_X1 port map( A1 => n14813, A2 => n11168, ZN => n11169);
   U4442 : AOI22_X1 port map( A1 => n11172, A2 => n11171, B1 => n10974, B2 => 
                           n11786, ZN => n11188);
   U4443 : XNOR2_X1 port map( A => n11174, B => n11173, ZN => n11177);
   U4444 : INV_X1 port map( A => n11175, ZN => n11176);
   U4445 : XNOR2_X1 port map( A => n11177, B => n11176, ZN => n11187);
   U4446 : NAND2_X1 port map( A1 => n11188, A2 => n11187, ZN => n11812);
   U4447 : MUX2_X1 port map( A => n14728, B => n13980, S => n12764, Z => n11180
                           );
   U4448 : XNOR2_X1 port map( A => n11272, B => n12014, ZN => n11178);
   U4449 : NAND2_X1 port map( A1 => n11178, A2 => n14786, ZN => n11179);
   U4450 : NAND2_X1 port map( A1 => n11180, A2 => n11179, ZN => n11185);
   U4451 : MUX2_X1 port map( A => n10940, B => n14020, S => n10869, Z => n11182
                           );
   U4452 : NAND2_X1 port map( A1 => n12230, A2 => n14477, ZN => n11181);
   U4453 : NAND2_X1 port map( A1 => n11182, A2 => n11181, ZN => n11186);
   U4454 : MUX2_X1 port map( A => n13449, B => n13448, S => n13914, Z => n11184
                           );
   U4455 : MUX2_X1 port map( A => n14833, B => n13451, S => n14785, Z => n11183
                           );
   U4456 : NAND2_X1 port map( A1 => n11184, A2 => n11183, ZN => n11789);
   U4457 : NAND2_X1 port map( A1 => n11812, A2 => n11813, ZN => n11189);
   U4458 : NAND2_X1 port map( A1 => n11189, A2 => n11811, ZN => n11433);
   U4459 : NAND2_X1 port map( A1 => n11431, A2 => n11433, ZN => n11193);
   U4460 : NAND2_X1 port map( A1 => n11193, A2 => n11432, ZN => n13898);
   U4461 : MUX2_X1 port map( A => n13449, B => n13448, S => n10904, Z => n11195
                           );
   U4462 : MUX2_X1 port map( A => n14833, B => n12783, S => n13924, Z => n11194
                           );
   U4463 : NAND2_X1 port map( A1 => n11195, A2 => n11194, ZN => n11200);
   U4464 : MUX2_X1 port map( A => n10640, B => n13868, S => n14819, Z => n11198
                           );
   U4465 : XNOR2_X1 port map( A => n12010, B => n12764, ZN => n11196);
   U4466 : NAND2_X1 port map( A1 => n14813, A2 => n11196, ZN => n11197);
   U4467 : NAND2_X1 port map( A1 => n11198, A2 => n11197, ZN => n11199);
   U4468 : NAND2_X1 port map( A1 => n11200, A2 => n11199, ZN => n11330);
   U4469 : NAND2_X1 port map( A1 => n11332, A2 => n11330, ZN => n11204);
   U4470 : BUF_X1 port map( A => n8332, Z => n13364);
   U4471 : MUX2_X1 port map( A => n14017, B => n13984, S => n13364, Z => n11203
                           );
   U4472 : MUX2_X1 port map( A => n14779, B => n14456, S => n14945, Z => n11202
                           );
   U4473 : AND2_X1 port map( A1 => n11203, A2 => n11202, ZN => n11329);
   U4474 : XNOR2_X1 port map( A => n11204, B => n11329, ZN => n11212);
   U4475 : NAND2_X1 port map( A1 => n14114, A2 => n10864, ZN => n11205);
   U4476 : NAND2_X1 port map( A1 => n11205, A2 => n10713, ZN => n11336);
   U4477 : MUX2_X1 port map( A => n14020, B => n14021, S => n13239, Z => n11207
                           );
   U4478 : NAND2_X1 port map( A1 => n14771, A2 => n10831, ZN => n11206);
   U4479 : NAND2_X1 port map( A1 => n11207, A2 => n11206, ZN => n11335);
   U4480 : XNOR2_X1 port map( A => n11336, B => n10677, ZN => n11210);
   U4481 : MUX2_X1 port map( A => n13362, B => n14114, S => n14594, Z => n11338
                           );
   U4482 : MUX2_X1 port map( A => n12146, B => n11225, S => n14719, Z => n11208
                           );
   U4483 : NOR2_X1 port map( A1 => n11338, A2 => n11208, ZN => n11209);
   U4484 : XNOR2_X1 port map( A => n11210, B => n11209, ZN => n11211);
   U4485 : NAND2_X1 port map( A1 => n11212, A2 => n11211, ZN => n11357);
   U4486 : NAND2_X1 port map( A1 => n11357, A2 => n11355, ZN => n11218);
   U4487 : NAND2_X1 port map( A1 => n11214, A2 => n11213, ZN => n11217);
   U4488 : NAND2_X1 port map( A1 => n11217, A2 => n11216, ZN => n11356);
   U4489 : XNOR2_X1 port map( A => n11218, B => n11356, ZN => n13897);
   U4490 : XNOR2_X1 port map( A => n13898, B => n13897, ZN => n11219);
   U4491 : XNOR2_X1 port map( A => n10678, B => n11219, ZN => n11483);
   U4492 : MUX2_X1 port map( A => n13371, B => n13372, S => n10869, Z => n11221
                           );
   U4493 : MUX2_X1 port map( A => n10641, B => n13373, S => n14477, Z => n11220
                           );
   U4494 : NAND2_X1 port map( A1 => n11221, A2 => n11220, ZN => n11261);
   U4495 : INV_X1 port map( A => n11261, ZN => n11233);
   U4496 : MUX2_X1 port map( A => n14833, B => n12783, S => n13810, Z => n11224
                           );
   U4497 : NAND2_X1 port map( A1 => n11222, A2 => n14727, ZN => n11223);
   U4498 : NAND2_X1 port map( A1 => n11224, A2 => n11223, ZN => n11259);
   U4499 : MUX2_X1 port map( A => n10713, B => n10636, S => n13273, Z => n11229
                           );
   U4500 : XOR2_X1 port map( A => n11226, B => n10913, Z => n11227);
   U4501 : NAND2_X1 port map( A1 => n11227, A2 => n14479, ZN => n11228);
   U4502 : NAND2_X1 port map( A1 => n11229, A2 => n11228, ZN => n11260);
   U4503 : NAND2_X1 port map( A1 => n11259, A2 => n11260, ZN => n11232);
   U4504 : INV_X1 port map( A => n11259, ZN => n11231);
   U4505 : INV_X1 port map( A => n11260, ZN => n11230);
   U4506 : AOI22_X1 port map( A1 => n11233, A2 => n11232, B1 => n11231, B2 => 
                           n11230, ZN => n11243);
   U4507 : MUX2_X1 port map( A => n10725, B => n11834, S => n8334, Z => n11236)
                           ;
   U4508 : XNOR2_X1 port map( A => n14117, B => n10861, ZN => n11234);
   U4509 : NAND2_X1 port map( A1 => n10857, A2 => n11234, ZN => n11235);
   U4510 : NAND2_X1 port map( A1 => n11236, A2 => n11235, ZN => n11263);
   U4511 : NAND2_X1 port map( A1 => n10635, A2 => n13809, ZN => n11262);
   U4512 : AND2_X1 port map( A1 => n11263, A2 => n11262, ZN => n11240);
   U4513 : NAND2_X1 port map( A1 => n10697, A2 => n11861, ZN => n11650);
   U4514 : NAND2_X1 port map( A1 => n10697, A2 => n14463, ZN => n11343);
   U4515 : BUF_X2 port map( A => n11343, Z => n13346);
   U4516 : MUX2_X1 port map( A => n12805, B => n13346, S => n10831, Z => n11239
                           );
   U4517 : MUX2_X1 port map( A => n13283, B => n14716, S => n12246, Z => n11238
                           );
   U4518 : NAND2_X1 port map( A1 => n11239, A2 => n11238, ZN => n11264);
   U4519 : OAI22_X1 port map( A1 => n11240, A2 => n11264, B1 => n11262, B2 => 
                           n11263, ZN => n11242);
   U4520 : INV_X1 port map( A => n11242, ZN => n11241);
   U4521 : NAND2_X1 port map( A1 => n10688, A2 => n11241, ZN => n11669);
   U4522 : NAND2_X1 port map( A1 => n11669, A2 => n11670, ZN => n11258);
   U4523 : MUX2_X1 port map( A => n14840, B => n10645, S => n8351, Z => n11244)
                           ;
   U4524 : NOR2_X1 port map( A1 => n11244, A2 => n14121, ZN => n11246);
   U4525 : INV_X1 port map( A => n10737, ZN => n12243);
   U4526 : INV_X1 port map( A => n13442, ZN => n11513);
   U4527 : MUX2_X1 port map( A => n12243, B => n11513, S => n11738, Z => n11245
                           );
   U4528 : NOR2_X1 port map( A1 => n11246, A2 => n11245, ZN => n11250);
   U4529 : MUX2_X1 port map( A => n8363, B => n10841, S => n12014, Z => n11247)
                           ;
   U4530 : INV_X1 port map( A => n11096, ZN => n11249);
   U4531 : NAND2_X1 port map( A1 => n11250, A2 => n11251, ZN => n11267);
   U4532 : INV_X1 port map( A => n11250, ZN => n11253);
   U4533 : NAND2_X1 port map( A1 => n11253, A2 => n11252, ZN => n11266);
   U4534 : MUX2_X1 port map( A => n12163, B => n14878, S => n10904, Z => n11254
                           );
   U4535 : NAND2_X1 port map( A1 => n11255, A2 => n11254, ZN => n11268);
   U4536 : INV_X1 port map( A => n11268, ZN => n11256);
   U4537 : NAND2_X1 port map( A1 => n11266, A2 => n11256, ZN => n11257);
   U4538 : NAND2_X1 port map( A1 => n11267, A2 => n11257, ZN => n11668);
   U4539 : XNOR2_X1 port map( A => n11258, B => n11668, ZN => n13209);
   U4540 : XNOR2_X1 port map( A => n11263, B => n11262, ZN => n11265);
   U4541 : XNOR2_X1 port map( A => n11264, B => n11265, ZN => n11269);
   U4542 : NAND2_X1 port map( A1 => n13563, A2 => n10888, ZN => n11270);
   U4543 : NAND2_X1 port map( A1 => n11270, A2 => n13562, ZN => n13210);
   U4544 : MUX2_X1 port map( A => n14840, B => n14118, S => n13273, Z => n11271
                           );
   U4545 : NOR2_X1 port map( A1 => n11271, A2 => n14121, ZN => n11274);
   U4546 : INV_X1 port map( A => n11282, ZN => n11278);
   U4547 : INV_X1 port map( A => n10680, ZN => n11275);
   U4548 : MUX2_X1 port map( A => n11275, B => n10638, S => n10841, Z => n11280
                           );
   U4549 : MUX2_X1 port map( A => n10725, B => n11834, S => n14117, Z => n11276
                           );
   U4550 : INV_X1 port map( A => n11276, ZN => n11279);
   U4551 : OR2_X1 port map( A1 => n11280, A2 => n11279, ZN => n11277);
   U4552 : NAND2_X1 port map( A1 => n11278, A2 => n11277, ZN => n13495);
   U4553 : NOR2_X1 port map( A1 => n11280, A2 => n11279, ZN => n11281);
   U4554 : NAND2_X1 port map( A1 => n11282, A2 => n11281, ZN => n13497);
   U4555 : NAND2_X1 port map( A1 => n13495, A2 => n13497, ZN => n11286);
   U4556 : MUX2_X1 port map( A => n13824, B => n12163, S => n14819, Z => n11284
                           );
   U4557 : NAND2_X1 port map( A1 => n11285, A2 => n11284, ZN => n13493);
   U4558 : XNOR2_X1 port map( A => n11286, B => n13493, ZN => n13499);
   U4559 : MUX2_X1 port map( A => n13346, B => n12805, S => n13813, Z => n13481
                           );
   U4560 : MUX2_X1 port map( A => n13347, B => n14716, S => n14478, Z => n13480
                           );
   U4561 : NAND2_X1 port map( A1 => n13481, A2 => n13480, ZN => n11289);
   U4562 : XNOR2_X1 port map( A => n8401, B => n13914, ZN => n11287);
   U4563 : NOR2_X1 port map( A1 => n11287, A2 => n13482, ZN => n11288);
   U4564 : XNOR2_X1 port map( A => n11289, B => n11288, ZN => n13500);
   U4565 : XNOR2_X1 port map( A => n13499, B => n13500, ZN => n11296);
   U4566 : MUX2_X1 port map( A => n10633, B => n10630, S => n10742, Z => n11291
                           );
   U4567 : MUX2_X1 port map( A => n10713, B => n10636, S => n10913, Z => n11290
                           );
   U4568 : NAND2_X1 port map( A1 => n11291, A2 => n11290, ZN => n13510);
   U4569 : XOR2_X1 port map( A => n13968, B => n13510, Z => n11294);
   U4570 : INV_X1 port map( A => FP_B(19), ZN => n10842);
   U4571 : MUX2_X1 port map( A => n13449, B => n13448, S => n10631, Z => n11293
                           );
   U4572 : MUX2_X1 port map( A => n14833, B => n12783, S => n8329, Z => n11292)
                           ;
   U4573 : NAND2_X1 port map( A1 => n11293, A2 => n11292, ZN => n13509);
   U4574 : XNOR2_X1 port map( A => n11294, B => n13509, ZN => n13501);
   U4575 : INV_X1 port map( A => n13501, ZN => n11295);
   U4576 : XNOR2_X1 port map( A => n11296, B => n11295, ZN => n13212);
   U4577 : OAI21_X1 port map( B1 => n13209, B2 => n13210, A => n13212, ZN => 
                           n11298);
   U4578 : NAND2_X1 port map( A1 => n13209, A2 => n13210, ZN => n11297);
   U4579 : NAND2_X1 port map( A1 => n11298, A2 => n11297, ZN => n11676);
   U4580 : NAND2_X1 port map( A1 => n14894, A2 => n14893, ZN => n12253);
   U4581 : NOR2_X1 port map( A1 => n12252, A2 => n14896, ZN => n12095);
   U4582 : NAND2_X1 port map( A1 => n10942, A2 => n12095, ZN => n14328);
   U4583 : OAI211_X1 port map( C1 => n8371, C2 => n10975, A => n8381, B => 
                           n14471, ZN => n11299);
   U4584 : MUX2_X1 port map( A => n14512, B => n8371, S => n10975, Z => n12249)
                           ;
   U4585 : NAND2_X1 port map( A1 => n12250, A2 => n12249, ZN => n12248);
   U4586 : MUX2_X1 port map( A => n8374, B => n2602, S => SIG_in_27_port, Z => 
                           n14331);
   U4587 : OR2_X1 port map( A1 => n12248, A2 => n14331, ZN => n12098);
   U4588 : MUX2_X1 port map( A => n14520, B => n2602, S => n10975, Z => n12097)
                           ;
   U4589 : OR2_X2 port map( A1 => n12098, A2 => n12097, ZN => n14338);
   U4590 : MUX2_X1 port map( A => n8345, B => n14497, S => SIG_in_27_port, Z =>
                           n14340);
   U4591 : MUX2_X1 port map( A => n14497, B => n8346, S => SIG_in_27_port, Z =>
                           n14339);
   U4592 : NAND2_X1 port map( A1 => n14340, A2 => n14339, ZN => n11300);
   U4593 : NOR2_X2 port map( A1 => n14338, A2 => n11300, ZN => n14345);
   U4594 : MUX2_X1 port map( A => n14513, B => n8346, S => n10975, Z => n14343)
                           ;
   U4595 : NAND2_X1 port map( A1 => n14345, A2 => n14343, ZN => n12194);
   U4596 : MUX2_X1 port map( A => n2598, B => n2597, S => n14730, Z => n12193);
   U4597 : OR2_X2 port map( A1 => n12194, A2 => n12193, ZN => n14346);
   U4598 : MUX2_X1 port map( A => n14515, B => n8391, S => n14730, Z => n14347)
                           ;
   U4599 : MUX2_X1 port map( A => n2597, B => n2596, S => n14730, Z => n11301);
   U4600 : INV_X1 port map( A => n11301, ZN => n14348);
   U4601 : NAND2_X1 port map( A1 => n14347, A2 => n14348, ZN => n11302);
   U4602 : NOR2_X2 port map( A1 => n14346, A2 => n11302, ZN => n14353);
   U4603 : MUX2_X1 port map( A => n14514, B => n8391, S => n10975, Z => n14351)
                           ;
   U4604 : NAND2_X1 port map( A1 => n14353, A2 => n14351, ZN => n14355);
   U4605 : MUX2_X1 port map( A => n2594, B => n2593, S => n14729, Z => n14354);
   U4607 : NAND2_X1 port map( A1 => n14457, A2 => n14818, ZN => n11303);
   U4608 : NAND2_X1 port map( A1 => n11304, A2 => n11303, ZN => n11495);
   U4609 : NAND2_X1 port map( A1 => n10857, A2 => n14738, ZN => n11494);
   U4610 : NAND2_X1 port map( A1 => n11495, A2 => n11494, ZN => n11493);
   U4611 : OR2_X1 port map( A1 => n14709, A2 => n2638, ZN => n10863);
   U4612 : INV_X1 port map( A => n11492, ZN => n11497);
   U4613 : XNOR2_X1 port map( A => n11493, B => n11497, ZN => n11311);
   U4614 : NAND2_X1 port map( A1 => n14739, A2 => n14731, ZN => n11306);
   U4615 : NAND2_X1 port map( A1 => n11306, A2 => n14725, ZN => n11310);
   U4616 : NAND2_X1 port map( A1 => n14741, A2 => n14448, ZN => n11307);
   U4617 : NAND2_X1 port map( A1 => n11307, A2 => n12018, ZN => n11309);
   U4618 : XNOR2_X1 port map( A => n8352, B => n11861, ZN => n11308);
   U4619 : AOI22_X1 port map( A1 => n11310, A2 => n11309, B1 => n12174, B2 => 
                           n11308, ZN => n11498);
   U4620 : XNOR2_X1 port map( A => n11311, B => n11498, ZN => n11328);
   U4621 : NAND2_X1 port map( A1 => n14482, A2 => n14771, ZN => n11315);
   U4622 : NAND2_X1 port map( A1 => n11313, A2 => n11312, ZN => n11314);
   U4623 : NAND2_X1 port map( A1 => n11315, A2 => n11314, ZN => n11500);
   U4624 : NAND2_X1 port map( A1 => n10641, A2 => n14785, ZN => n11317);
   U4625 : NAND2_X1 port map( A1 => n12639, A2 => n14593, ZN => n11316);
   U4626 : NAND2_X1 port map( A1 => n11317, A2 => n11316, ZN => n11320);
   U4627 : XNOR2_X1 port map( A => n8350, B => n14713, ZN => n11318);
   U4628 : NAND2_X1 port map( A1 => n11318, A2 => n12640, ZN => n11319);
   U4629 : NAND2_X1 port map( A1 => n11320, A2 => n11319, ZN => n11501);
   U4630 : XNOR2_X1 port map( A => n11501, B => n11500, ZN => n11326);
   U4631 : MUX2_X1 port map( A => n12146, B => n11225, S => n14777, Z => n11324
                           );
   U4632 : XNOR2_X1 port map( A => n11321, B => n14447, ZN => n11322);
   U4633 : INV_X1 port map( A => n11504, ZN => n11325);
   U4634 : XNOR2_X1 port map( A => n11326, B => n11325, ZN => n11327);
   U4635 : NAND2_X1 port map( A1 => n11328, A2 => n11327, ZN => n11562);
   U4636 : NAND2_X1 port map( A1 => n11563, A2 => n11562, ZN => n11352);
   U4637 : NAND2_X1 port map( A1 => n11330, A2 => n11329, ZN => n11331);
   U4638 : NAND2_X1 port map( A1 => n11332, A2 => n11331, ZN => n11561);
   U4639 : XNOR2_X1 port map( A => n10723, B => n11561, ZN => n11350);
   U4640 : NAND2_X1 port map( A1 => n11336, A2 => n11335, ZN => n11334);
   U4641 : AOI22_X1 port map( A1 => n11225, A2 => n14719, B1 => n12146, B2 => 
                           n10864, ZN => n11333);
   U4642 : NAND2_X1 port map( A1 => n11334, A2 => n11333, ZN => n11339);
   U4643 : OAI21_X1 port map( B1 => n11339, B2 => n11338, A => n11337, ZN => 
                           n11559);
   U4644 : MUX2_X1 port map( A => n11096, B => n13908, S => n14449, Z => n11342
                           );
   U4645 : MUX2_X1 port map( A => n13920, B => n14728, S => n14477, Z => n11340
                           );
   U4646 : INV_X1 port map( A => n11340, ZN => n11341);
   U4647 : OR2_X1 port map( A1 => n11342, A2 => n11341, ZN => n11556);
   U4648 : XNOR2_X1 port map( A => n11559, B => n11556, ZN => n11348);
   U4649 : NAND2_X1 port map( A1 => n11345, A2 => n11344, ZN => n11405);
   U4650 : MUX2_X1 port map( A => n11043, B => n11957, S => n11965, Z => n11347
                           );
   U4651 : MUX2_X1 port map( A => n10725, B => n11149, S => n11272, Z => n11346
                           );
   U4652 : NAND2_X1 port map( A1 => n11347, A2 => n11346, ZN => n13885);
   U4653 : INV_X1 port map( A => n11555, ZN => n11557);
   U4654 : XNOR2_X1 port map( A => n11557, B => n11348, ZN => n11353);
   U4655 : INV_X1 port map( A => n11353, ZN => n11349);
   U4656 : NAND2_X1 port map( A1 => n11350, A2 => n11349, ZN => n12261);
   U4657 : INV_X1 port map( A => n11561, ZN => n11351);
   U4658 : XNOR2_X1 port map( A => n11352, B => n11351, ZN => n11354);
   U4659 : NAND2_X1 port map( A1 => n11354, A2 => n11353, ZN => n12259);
   U4660 : NAND2_X1 port map( A1 => n12261, A2 => n12259, ZN => n11359);
   U4661 : NAND2_X1 port map( A1 => n11356, A2 => n11355, ZN => n11358);
   U4662 : NAND2_X1 port map( A1 => n11358, A2 => n11357, ZN => n12260);
   U4663 : MUX2_X1 port map( A => n13283, B => n14716, S => n14785, Z => n11362
                           );
   U4664 : NAND2_X1 port map( A1 => n14479, A2 => n14719, ZN => n13881);
   U4665 : MUX2_X1 port map( A => n11043, B => n10680, S => n8351, Z => n11361)
                           ;
   U4666 : MUX2_X1 port map( A => n10725, B => n11834, S => n12764, Z => n11360
                           );
   U4667 : AND2_X1 port map( A1 => n11361, A2 => n11360, ZN => n13882);
   U4668 : INV_X1 port map( A => n11362, ZN => n11364);
   U4669 : INV_X1 port map( A => n13881, ZN => n11363);
   U4670 : NAND2_X1 port map( A1 => n11364, A2 => n11363, ZN => n11365);
   U4671 : OAI211_X1 port map( C1 => n11366, C2 => n13881, A => n13882, B => 
                           n11365, ZN => n11367);
   U4672 : NAND2_X1 port map( A1 => n11368, A2 => n11367, ZN => n13186);
   U4673 : AOI21_X1 port map( B1 => n14832, B2 => n14448, A => n13265, ZN => 
                           n11374);
   U4674 : NAND2_X1 port map( A1 => FP_B(5), A2 => FP_A(10), ZN => n10852);
   U4675 : OAI21_X1 port map( B1 => n11369, B2 => n14725, A => n12124, ZN => 
                           n11370);
   U4676 : INV_X1 port map( A => n11370, ZN => n11373);
   U4677 : NAND2_X1 port map( A1 => n11371, A2 => n14727, ZN => n11372);
   U4678 : OAI21_X1 port map( B1 => n11374, B2 => n11373, A => n11372, ZN => 
                           n13877);
   U4679 : MUX2_X1 port map( A => n14021, B => n14020, S => n10831, Z => n11376
                           );
   U4680 : NAND2_X1 port map( A1 => n14452, A2 => n12230, ZN => n11375);
   U4681 : NAND2_X1 port map( A1 => n11376, A2 => n11375, ZN => n13878);
   U4682 : MUX2_X1 port map( A => n10745, B => n12142, S => n14594, Z => n11379
                           );
   U4683 : XNOR2_X1 port map( A => n14447, B => n12671, ZN => n11377);
   U4684 : NAND2_X1 port map( A1 => n12640, A2 => n11377, ZN => n11378);
   U4685 : AND2_X1 port map( A1 => n11379, A2 => n11378, ZN => n13879);
   U4686 : INV_X1 port map( A => n13877, ZN => n11382);
   U4687 : INV_X1 port map( A => n13878, ZN => n11381);
   U4688 : NAND2_X1 port map( A1 => n11382, A2 => n11381, ZN => n11383);
   U4689 : NAND2_X1 port map( A1 => n11384, A2 => n11383, ZN => n13184);
   U4690 : NAND2_X1 port map( A1 => n13868, A2 => n14451, ZN => n11387);
   U4691 : NAND2_X1 port map( A1 => n10640, A2 => n10904, ZN => n11386);
   U4692 : NAND2_X1 port map( A1 => n11387, A2 => n11386, ZN => n11391);
   U4693 : XOR2_X1 port map( A => B_SIG_8_port, B => n12124, Z => n11389);
   U4694 : NAND2_X1 port map( A1 => n14813, A2 => n11389, ZN => n11390);
   U4695 : NAND2_X1 port map( A1 => n11391, A2 => n11390, ZN => n13873);
   U4696 : MUX2_X1 port map( A => n14728, B => n13980, S => n11965, Z => n11394
                           );
   U4697 : XNOR2_X1 port map( A => n10913, B => n12014, ZN => n11392);
   U4698 : NAND2_X1 port map( A1 => n14786, A2 => n11392, ZN => n11393);
   U4699 : NAND2_X1 port map( A1 => n11394, A2 => n11393, ZN => n13872);
   U4700 : AND2_X1 port map( A1 => n13872, A2 => n13873, ZN => n11397);
   U4701 : MUX2_X1 port map( A => n11201, B => n14017, S => n10869, Z => n11396
                           );
   U4702 : MUX2_X1 port map( A => n13915, B => n14779, S => n10742, Z => n11395
                           );
   U4703 : NAND2_X1 port map( A1 => n11396, A2 => n11395, ZN => n13874);
   U4704 : OAI22_X1 port map( A1 => n11397, A2 => n13874, B1 => n13873, B2 => 
                           n13872, ZN => n13183);
   U4705 : OAI21_X1 port map( B1 => n13186, B2 => n13184, A => n13183, ZN => 
                           n11399);
   U4706 : NAND2_X1 port map( A1 => n13186, A2 => n13184, ZN => n11398);
   U4707 : NAND2_X1 port map( A1 => n11399, A2 => n11398, ZN => n11546);
   U4708 : MUX2_X1 port map( A => n13371, B => n13372, S => n14593, Z => n11401
                           );
   U4709 : MUX2_X1 port map( A => n10745, B => n13373, S => n14025, Z => n11400
                           );
   U4710 : NAND2_X1 port map( A1 => n11401, A2 => n11400, ZN => n13888);
   U4711 : MUX2_X1 port map( A => n13920, B => n14728, S => n14455, Z => n11404
                           );
   U4712 : XNOR2_X1 port map( A => n10742, B => n12014, ZN => n11402);
   U4713 : NAND2_X1 port map( A1 => n14786, A2 => n11402, ZN => n11403);
   U4714 : NAND2_X1 port map( A1 => n11404, A2 => n11403, ZN => n11409);
   U4715 : AND2_X1 port map( A1 => n13888, A2 => n11409, ZN => n11413);
   U4716 : INV_X1 port map( A => n13884, ZN => n11408);
   U4717 : NAND2_X1 port map( A1 => n13888, A2 => n11409, ZN => n11407);
   U4718 : NAND3_X1 port map( A1 => n11408, A2 => n11407, A3 => n11406, ZN => 
                           n11412);
   U4719 : INV_X1 port map( A => n13888, ZN => n11410);
   U4720 : INV_X1 port map( A => n11409, ZN => n13887);
   U4721 : NAND2_X1 port map( A1 => n11410, A2 => n13887, ZN => n11411);
   U4722 : OAI211_X1 port map( C1 => n11413, C2 => n11557, A => n11412, B => 
                           n11411, ZN => n11414);
   U4723 : INV_X1 port map( A => n11414, ZN => n11427);
   U4724 : MUX2_X1 port map( A => n10640, B => n13868, S => n14453, Z => n11417
                           );
   U4725 : INV_X1 port map( A => n14464, ZN => n13328);
   U4726 : XNOR2_X1 port map( A => n12010, B => n13328, ZN => n11415);
   U4727 : NAND2_X1 port map( A1 => n14813, A2 => n11415, ZN => n11416);
   U4728 : MUX2_X1 port map( A => n11201, B => n14017, S => n10831, Z => n11420
                           );
   U4729 : MUX2_X1 port map( A => n13915, B => n14779, S => n13364, Z => n11419
                           );
   U4730 : XNOR2_X1 port map( A => n11526, B => n11524, ZN => n11425);
   U4731 : MUX2_X1 port map( A => n14833, B => n12783, S => n13485, Z => n11421
                           );
   U4732 : XOR2_X1 port map( A => B_SIG_8_port, B => n14725, Z => n11422);
   U4733 : INV_X1 port map( A => n11528, ZN => n11424);
   U4734 : XNOR2_X1 port map( A => n11425, B => n11424, ZN => n11426);
   U4735 : NAND2_X1 port map( A1 => n11427, A2 => n11426, ZN => n11545);
   U4736 : NAND2_X1 port map( A1 => n11545, A2 => n11544, ZN => n11428);
   U4737 : XNOR2_X1 port map( A => n11546, B => n11428, ZN => n12042);
   U4738 : XNOR2_X1 port map( A => intadd_66_n2, B => n12042, ZN => n11429);
   U4739 : XNOR2_X1 port map( A => n10744, B => n11429, ZN => 
                           intadd_66_SUM_2_port);
   U4743 : NOR2_X1 port map( A1 => n12342, A2 => n14684, ZN => n11430);
   U4744 : INV_X1 port map( A => n11430, ZN => n12046);
   U4745 : NAND2_X1 port map( A1 => n11432, A2 => n11431, ZN => n11434);
   U4746 : XNOR2_X1 port map( A => n11434, B => n11433, ZN => n13195);
   U4747 : NAND2_X1 port map( A1 => n11436, A2 => n11435, ZN => n11439);
   U4748 : INV_X1 port map( A => n11437, ZN => n11438);
   U4749 : XNOR2_X1 port map( A => n11439, B => n11438, ZN => n11479);
   U4750 : INV_X1 port map( A => n11440, ZN => n11445);
   U4751 : NAND2_X1 port map( A1 => n11462, A2 => n11441, ZN => n11443);
   U4752 : NAND2_X1 port map( A1 => n11443, A2 => n11442, ZN => n11444);
   U4753 : XNOR2_X1 port map( A => n11445, B => n11444, ZN => n11448);
   U4754 : INV_X1 port map( A => n11446, ZN => n11447);
   U4755 : XNOR2_X1 port map( A => n11448, B => n11447, ZN => n11478);
   U4756 : NAND2_X1 port map( A1 => n11479, A2 => n11478, ZN => n11816);
   U4757 : MUX2_X1 port map( A => n13347, B => n14716, S => n14719, Z => n11451
                           );
   U4758 : XNOR2_X1 port map( A => n14463, B => n14594, ZN => n11449);
   U4759 : NAND2_X1 port map( A1 => n12174, A2 => n11449, ZN => n11450);
   U4760 : MUX2_X1 port map( A => n14833, B => n12783, S => n14447, Z => n11454
                           );
   U4761 : XNOR2_X1 port map( A => n14725, B => n14593, ZN => n11452);
   U4762 : NAND2_X1 port map( A1 => n14727, A2 => n11452, ZN => n11453);
   U4763 : NAND2_X1 port map( A1 => n11454, A2 => n11453, ZN => n11721);
   U4764 : MUX2_X1 port map( A => n14020, B => n10939, S => n10742, Z => n11456
                           );
   U4765 : NAND2_X1 port map( A1 => n14771, A2 => n14455, ZN => n11455);
   U4766 : NAND2_X1 port map( A1 => n11456, A2 => n11455, ZN => n11457);
   U4767 : NAND2_X1 port map( A1 => n11721, A2 => n11457, ZN => n11459);
   U4768 : INV_X1 port map( A => n11721, ZN => n11458);
   U4769 : XNOR2_X1 port map( A => n11461, B => n11460, ZN => n11463);
   U4770 : XNOR2_X1 port map( A => n11463, B => n11462, ZN => n11475);
   U4771 : MUX2_X1 port map( A => n11096, B => n13908, S => n11738, Z => n11466
                           );
   U4772 : MUX2_X1 port map( A => n13920, B => n14728, S => n14819, Z => n11464
                           );
   U4773 : INV_X1 port map( A => n11464, ZN => n11465);
   U4774 : OR2_X1 port map( A1 => n11466, A2 => n11465, ZN => n11690);
   U4775 : XOR2_X1 port map( A => n12124, B => n14731, Z => n11467);
   U4776 : NAND2_X1 port map( A1 => n11467, A2 => n14813, ZN => n11469);
   U4777 : MUX2_X1 port map( A => n10640, B => n13868, S => n14465, Z => n11468
                           );
   U4778 : NAND2_X1 port map( A1 => n11469, A2 => n11468, ZN => n11473);
   U4779 : MUX2_X1 port map( A => n14017, B => n11201, S => n12743, Z => n11471
                           );
   U4780 : MUX2_X1 port map( A => n13915, B => n14779, S => n8351, Z => n11470)
                           ;
   U4781 : NAND2_X1 port map( A1 => n11471, A2 => n11470, ZN => n11472);
   U4782 : OAI21_X1 port map( B1 => n11690, B2 => n11474, A => n11692, ZN => 
                           n11802);
   U4783 : NAND2_X1 port map( A1 => n11800, A2 => n11802, ZN => n11477);
   U4784 : NAND2_X1 port map( A1 => n11477, A2 => n11801, ZN => n13891);
   U4785 : NAND2_X1 port map( A1 => n11816, A2 => n13891, ZN => n11480);
   U4786 : OR2_X1 port map( A1 => n11479, A2 => n11478, ZN => n11817);
   U4787 : NAND2_X1 port map( A1 => n11480, A2 => n11817, ZN => n13196);
   U4788 : OAI21_X1 port map( B1 => n13195, B2 => n13196, A => 
                           intadd_56_A_3_port, ZN => n11482);
   U4789 : NAND2_X1 port map( A1 => n13195, A2 => n13196, ZN => n11481);
   U4790 : NAND2_X1 port map( A1 => n10750, A2 => n10748, ZN => n14753);
   U4791 : MUX2_X1 port map( A => n13347, B => n14716, S => n8352, Z => n11486)
                           ;
   U4792 : XNOR2_X1 port map( A => n13485, B => n10877, ZN => n11484);
   U4793 : NAND2_X1 port map( A1 => n11484, A2 => n12174, ZN => n11485);
   U4794 : NAND2_X1 port map( A1 => n11486, A2 => n11485, ZN => n11505);
   U4795 : AOI21_X1 port map( B1 => n10738, B2 => n14719, A => n14840, ZN => 
                           n11506);
   U4796 : NAND2_X1 port map( A1 => n11505, A2 => n11506, ZN => n13204);
   U4797 : MUX2_X1 port map( A => n14728, B => n13980, S => n13364, Z => n11490
                           );
   U4798 : XNOR2_X1 port map( A => FP_A(5), B => n360, ZN => n10830);
   U4799 : NAND2_X1 port map( A1 => n14786, A2 => n11488, ZN => n11489);
   U4800 : AND2_X1 port map( A1 => n11490, A2 => n11489, ZN => n13199);
   U4801 : XNOR2_X1 port map( A => n13204, B => n13199, ZN => n11491);
   U4802 : MUX2_X1 port map( A => n13372, B => n13371, S => n13924, Z => n13202
                           );
   U4803 : MUX2_X1 port map( A => n10745, B => n12142, S => n14448, Z => n13200
                           );
   U4804 : NAND2_X1 port map( A1 => n13202, A2 => n13200, ZN => n13206);
   U4805 : NAND2_X1 port map( A1 => n11493, A2 => n11492, ZN => n11499);
   U4806 : AND2_X1 port map( A1 => n11495, A2 => n11494, ZN => n11496);
   U4807 : NAND2_X1 port map( A1 => n11501, A2 => n11500, ZN => n11503);
   U4808 : NOR2_X1 port map( A1 => n11501, A2 => n11500, ZN => n11502);
   U4809 : AOI21_X1 port map( B1 => n11504, B2 => n11503, A => n11502, ZN => 
                           n11508);
   U4810 : NAND2_X1 port map( A1 => n11507, A2 => n11508, ZN => n11509);
   U4811 : OAI21_X1 port map( B1 => n11506, B2 => n11505, A => n13204, ZN => 
                           n11542);
   U4812 : INV_X1 port map( A => n11507, ZN => n11540);
   U4813 : INV_X1 port map( A => n11508, ZN => n11541);
   U4815 : XNOR2_X1 port map( A => n11511, B => n11512, ZN => n11518);
   U4816 : OAI22_X1 port map( A1 => n10864, A2 => n13442, B1 => n10738, B2 => 
                           n14719, ZN => n11516);
   U4817 : INV_X1 port map( A => n11514, ZN => n11515);
   U4818 : NOR2_X1 port map( A1 => n11516, A2 => n11515, ZN => n11517);
   U4819 : XNOR2_X1 port map( A => n11518, B => n11517, ZN => n11537);
   U4820 : INV_X1 port map( A => n11519, ZN => n11520);
   U4821 : XNOR2_X1 port map( A => n11521, B => n11520, ZN => n11523);
   U4822 : XNOR2_X1 port map( A => n11523, B => n11522, ZN => n11531);
   U4823 : NAND2_X1 port map( A1 => n11531, A2 => n11537, ZN => n11533);
   U4824 : INV_X1 port map( A => n11524, ZN => n11525);
   U4825 : OAI21_X1 port map( B1 => n11525, B2 => n11528, A => n11527, ZN => 
                           n11530);
   U4826 : NAND2_X1 port map( A1 => n11525, A2 => n11528, ZN => n11529);
   U4827 : NAND2_X1 port map( A1 => n11530, A2 => n11529, ZN => n11535);
   U4828 : INV_X1 port map( A => n11537, ZN => n11532);
   U4829 : INV_X1 port map( A => n11531, ZN => n11538);
   U4830 : AOI22_X1 port map( A1 => n11533, A2 => n11535, B1 => n11532, B2 => 
                           n11538, ZN => n13160);
   U4831 : INV_X1 port map( A => n13160, ZN => n11689);
   U4832 : XNOR2_X1 port map( A => n11689, B => n11534, ZN => n13623);
   U4833 : INV_X1 port map( A => n11535, ZN => n11536);
   U4834 : XNOR2_X1 port map( A => n11537, B => n11536, ZN => n11539);
   U4835 : XNOR2_X1 port map( A => n11539, B => n11538, ZN => n12960);
   U4836 : XNOR2_X1 port map( A => n11541, B => n11540, ZN => n11543);
   U4837 : OAI21_X1 port map( B1 => n10949, B2 => n11546, A => n11545, ZN => 
                           n12958);
   U4838 : INV_X1 port map( A => n10701, ZN => n11547);
   U4839 : OAI21_X1 port map( B1 => n12960, B2 => n12957, A => n11547, ZN => 
                           n13622);
   U4840 : NAND2_X1 port map( A1 => n12960, A2 => n12957, ZN => n13621);
   U4841 : INV_X1 port map( A => n11550, ZN => n11552);
   U4842 : NAND2_X1 port map( A1 => n11555, A2 => n11556, ZN => n11560);
   U4843 : INV_X1 port map( A => n11556, ZN => n11558);
   U4844 : AOI22_X1 port map( A1 => n11560, A2 => n11559, B1 => n11558, B2 => 
                           n11557, ZN => n11566);
   U4845 : NAND2_X1 port map( A1 => n11565, A2 => n11566, ZN => n12961);
   U4846 : NAND2_X1 port map( A1 => n11562, A2 => n11561, ZN => n11564);
   U4847 : NAND2_X1 port map( A1 => n11564, A2 => n11563, ZN => n12963);
   U4848 : NAND2_X1 port map( A1 => n12961, A2 => n12963, ZN => n11569);
   U4849 : INV_X1 port map( A => n11565, ZN => n11568);
   U4850 : INV_X1 port map( A => n11566, ZN => n11567);
   U4851 : NAND2_X1 port map( A1 => n11568, A2 => n11567, ZN => n12962);
   U4852 : XNOR2_X1 port map( A => n11570, B => n11678, ZN => n11575);
   U4853 : INV_X1 port map( A => n11571, ZN => n11572);
   U4854 : XNOR2_X1 port map( A => n11573, B => n11572, ZN => n11574);
   U4855 : XNOR2_X1 port map( A => n11574, B => intadd_46_SUM_0_port, ZN => 
                           n11683);
   U4857 : NAND2_X1 port map( A1 => n11578, A2 => n11577, ZN => n14769);
   U4858 : MUX2_X1 port map( A => n10633, B => n10630, S => n13273, Z => n11580
                           );
   U4859 : MUX2_X1 port map( A => n10713, B => n10636, S => n13328, Z => n11579
                           );
   U4860 : NAND2_X1 port map( A1 => n11580, A2 => n11579, ZN => n13063);
   U4861 : INV_X1 port map( A => n13063, ZN => n11590);
   U4862 : MUX2_X1 port map( A => n14833, B => n12783, S => n14478, Z => n11583
                           );
   U4863 : XNOR2_X1 port map( A => n12018, B => n13239, ZN => n11581);
   U4864 : NAND2_X1 port map( A1 => n11581, A2 => n14727, ZN => n11582);
   U4865 : NAND2_X1 port map( A1 => n11583, A2 => n11582, ZN => n13062);
   U4866 : MUX2_X1 port map( A => n13824, B => n12163, S => n14788, Z => n11586
                           );
   U4867 : XNOR2_X1 port map( A => n10905, B => n14715, ZN => n11584);
   U4868 : NAND2_X1 port map( A1 => n11584, A2 => n14789, ZN => n11585);
   U4869 : NAND2_X1 port map( A1 => n11586, A2 => n11585, ZN => n13061);
   U4870 : NAND2_X1 port map( A1 => n13062, A2 => n13061, ZN => n11589);
   U4871 : INV_X1 port map( A => n13062, ZN => n11588);
   U4872 : INV_X1 port map( A => n13061, ZN => n11587);
   U4873 : AOI22_X1 port map( A1 => n11590, A2 => n11589, B1 => n11588, B2 => 
                           n11587, ZN => n13571);
   U4874 : MUX2_X1 port map( A => n13372, B => n13371, S => n10742, Z => n11592
                           );
   U4875 : MUX2_X1 port map( A => n10641, B => n12142, S => n14455, Z => n11591
                           );
   U4876 : NAND2_X1 port map( A1 => n11592, A2 => n11591, ZN => n13059);
   U4877 : XOR2_X1 port map( A => n8334, B => n8355, Z => n11593);
   U4878 : NAND2_X1 port map( A1 => n11593, A2 => n10857, ZN => n11605);
   U4879 : MUX2_X1 port map( A => n10725, B => n11149, S => n13450, Z => n11606
                           );
   U4880 : NAND2_X1 port map( A1 => n11596, A2 => n11606, ZN => n13057);
   U4881 : NAND2_X1 port map( A1 => n13059, A2 => n13057, ZN => n11610);
   U4882 : XNOR2_X1 port map( A => n12124, B => n8325, ZN => n11601);
   U4883 : NOR2_X1 port map( A1 => n12125, A2 => A_SIG_8_port, ZN => n11597);
   U4884 : NAND3_X1 port map( A1 => n8355, A2 => n12125, A3 => A_SIG_8_port, ZN
                           => n11598);
   U4885 : AND2_X1 port map( A1 => n11598, A2 => n12010, ZN => n11599);
   U4886 : NAND2_X1 port map( A1 => n14017, A2 => n13915, ZN => n13054);
   U4887 : INV_X1 port map( A => n13054, ZN => n11608);
   U4888 : NAND2_X1 port map( A1 => n14728, A2 => n13920, ZN => n11603);
   U4889 : XNOR2_X1 port map( A => n12014, B => n14117, ZN => n12134);
   U4890 : XNOR2_X1 port map( A => n14881, B => n12014, ZN => n11602);
   U4891 : AOI22_X1 port map( A1 => n11603, A2 => n12134, B1 => n14786, B2 => 
                           n11602, ZN => n13055);
   U4892 : INV_X1 port map( A => n13055, ZN => n11604);
   U4893 : NAND2_X1 port map( A1 => n11613, A2 => n11604, ZN => n11609);
   U4894 : NAND2_X1 port map( A1 => n11606, A2 => n11605, ZN => n11607);
   U4895 : NAND2_X1 port map( A1 => n11607, A2 => n11594, ZN => n13058);
   U4896 : NAND2_X1 port map( A1 => n13571, A2 => n13569, ZN => n11616);
   U4897 : INV_X1 port map( A => n13059, ZN => n11611);
   U4898 : NAND2_X1 port map( A1 => n11611, A2 => n13058, ZN => n11615);
   U4899 : NAND2_X1 port map( A1 => n11612, A2 => n13055, ZN => n11614);
   U4900 : NAND4_X1 port map( A1 => n11615, A2 => n11614, A3 => n13057, A4 => 
                           n11613, ZN => n13570);
   U4901 : AND2_X1 port map( A1 => n11616, A2 => n13570, ZN => n11627);
   U4902 : INV_X1 port map( A => n11627, ZN => n11624);
   U4903 : MUX2_X1 port map( A => n13372, B => n13371, S => n13234, Z => n11618
                           );
   U4904 : MUX2_X1 port map( A => n10641, B => n13373, S => n14945, Z => n11617
                           );
   U4905 : NAND2_X1 port map( A1 => n11618, A2 => n11617, ZN => n13505);
   U4906 : BUF_X2 port map( A => n14880, Z => n13817);
   U4907 : MUX2_X1 port map( A => n13817, B => n10885, S => n10904, Z => n11620
                           );
   U4908 : NAND2_X1 port map( A1 => n14510, A2 => n14718, ZN => n11995);
   U4909 : BUF_X4 port map( A => n11995, Z => n13819);
   U4910 : MUX2_X1 port map( A => n13819, B => n14882, S => n13924, Z => n11619
                           );
   U4911 : NAND2_X1 port map( A1 => n11620, A2 => n11619, ZN => n13506);
   U4912 : XNOR2_X1 port map( A => n13505, B => n13506, ZN => n11625);
   U4913 : MUX2_X1 port map( A => n11743, B => n13323, S => n8334, Z => n11622)
                           ;
   U4915 : INV_X1 port map( A => n13868, ZN => n11933);
   U4916 : MUX2_X1 port map( A => n11385, B => n11933, S => n14458, Z => n11621
                           );
   U4917 : XOR2_X1 port map( A => n11625, B => n13504, Z => n11623);
   U4918 : NAND2_X1 port map( A1 => n11624, A2 => n11623, ZN => n13586);
   U4919 : XNOR2_X1 port map( A => n11625, B => n13504, ZN => n11626);
   U4920 : NAND2_X1 port map( A1 => n11627, A2 => n11626, ZN => n13585);
   U4921 : NAND2_X1 port map( A1 => n14716, A2 => n14449, ZN => n11630);
   U4922 : NAND2_X1 port map( A1 => n13283, A2 => n10869, ZN => n11629);
   U4923 : XNOR2_X1 port map( A => n13364, B => n10877, ZN => n11628);
   U4924 : AOI22_X1 port map( A1 => n11630, A2 => n11629, B1 => n11628, B2 => 
                           n12174, ZN => n11636);
   U4925 : NAND2_X1 port map( A1 => n14785, A2 => n13809, ZN => n11635);
   U4926 : NAND2_X1 port map( A1 => n11636, A2 => n11635, ZN => n12152);
   U4927 : NAND2_X1 port map( A1 => n13442, A2 => n11703, ZN => n11633);
   U4928 : NAND2_X1 port map( A1 => n10738, A2 => n14819, ZN => n11632);
   U4929 : XNOR2_X1 port map( A => n10693, B => n12764, ZN => n11631);
   U4930 : NAND2_X1 port map( A1 => n11637, A2 => n12151, ZN => n12188);
   U4931 : MUX2_X1 port map( A => n10640, B => n13868, S => n10726, Z => n11640
                           );
   U4932 : BUF_X2 port map( A => n8349, Z => n13450);
   U4933 : XNOR2_X1 port map( A => n12010, B => n13450, ZN => n11638);
   U4934 : NAND2_X1 port map( A1 => n14813, A2 => n11638, ZN => n11639);
   U4935 : NAND2_X1 port map( A1 => n11640, A2 => n11639, ZN => n11644);
   U4936 : MUX2_X1 port map( A => n13817, B => n10886, S => n8352, Z => n11642)
                           ;
   U4937 : MUX2_X1 port map( A => n11995, B => n14882, S => n14731, Z => n11641
                           );
   U4938 : NOR2_X1 port map( A1 => n11644, A2 => n11645, ZN => n12157);
   U4939 : INV_X1 port map( A => n12157, ZN => n11643);
   U4940 : NAND2_X1 port map( A1 => n12188, A2 => n11643, ZN => n11647);
   U4941 : INV_X1 port map( A => n12156, ZN => n11646);
   U4942 : NAND2_X1 port map( A1 => n11647, A2 => n11646, ZN => n13587);
   U4943 : INV_X1 port map( A => n11743, ZN => n13268);
   U4944 : INV_X1 port map( A => n13323, ZN => n11648);
   U4945 : MUX2_X1 port map( A => n13268, B => n11648, S => n13261, Z => n13432
                           );
   U4946 : MUX2_X1 port map( A => n10640, B => n13868, S => n14467, Z => n13431
                           );
   U4947 : NAND2_X1 port map( A1 => n13432, A2 => n13431, ZN => n13429);
   U4948 : MUX2_X1 port map( A => n13283, B => n14716, S => n13810, Z => n11654
                           );
   U4949 : INV_X1 port map( A => n11651, ZN => n11652);
   U4950 : MUX2_X1 port map( A => n12163, B => n14878, S => n12764, Z => n11655
                           );
   U4951 : NAND2_X1 port map( A1 => n11656, A2 => n11655, ZN => n13430);
   U4952 : XNOR2_X1 port map( A => n13433, B => n13430, ZN => n11657);
   U4953 : XNOR2_X1 port map( A => n11657, B => n13429, ZN => n11665);
   U4954 : MUX2_X1 port map( A => n13449, B => n13448, S => n13450, Z => n11659
                           );
   U4955 : MUX2_X1 port map( A => n14833, B => n12783, S => n13282, Z => n11658
                           );
   U4956 : NAND2_X1 port map( A1 => n11659, A2 => n11658, ZN => n13426);
   U4957 : MUX2_X1 port map( A => n13371, B => n13372, S => n10831, Z => n11661
                           );
   U4958 : MUX2_X1 port map( A => n13373, B => n10745, S => n13234, Z => n11660
                           );
   U4959 : NAND2_X1 port map( A1 => n11661, A2 => n11660, ZN => n13629);
   U4960 : MUX2_X1 port map( A => n10630, B => n10633, S => n10869, Z => n11663
                           );
   U4961 : MUX2_X1 port map( A => n10713, B => n10636, S => n10743, Z => n11662
                           );
   U4962 : NAND2_X1 port map( A1 => n11663, A2 => n11662, ZN => n13630);
   U4963 : NAND2_X1 port map( A1 => n11665, A2 => n11666, ZN => n13521);
   U4964 : INV_X1 port map( A => n11666, ZN => n11667);
   U4965 : NAND2_X1 port map( A1 => n10944, A2 => n11667, ZN => n13523);
   U4966 : NAND2_X1 port map( A1 => n13521, A2 => n13523, ZN => n11672);
   U4967 : NAND2_X1 port map( A1 => n11669, A2 => n11668, ZN => n11671);
   U4968 : NAND2_X1 port map( A1 => n11671, A2 => n11670, ZN => n13522);
   U4969 : XNOR2_X1 port map( A => n11672, B => n13522, ZN => n11673);
   U4970 : NAND2_X1 port map( A1 => n11674, A2 => n11673, ZN => n14254);
   U4971 : INV_X1 port map( A => n11674, ZN => n11675);
   U4972 : NAND2_X1 port map( A1 => n10945, A2 => n11675, ZN => n14253);
   U4973 : NAND2_X1 port map( A1 => n14254, A2 => n14253, ZN => n14199);
   U4974 : XNOR2_X1 port map( A => n14199, B => n11677, ZN => n14861);
   U4975 : NAND2_X1 port map( A1 => n14924, A2 => EXP_out_round_1_port, ZN => 
                           n14926);
   U4976 : XNOR2_X1 port map( A => n11680, B => n11679, ZN => n11681);
   U4977 : XNOR2_X1 port map( A => n11685, B => n11684, ZN => n12233);
   U4978 : AND2_X1 port map( A1 => n11686, A2 => n10894, ZN => n11687);
   U4979 : INV_X1 port map( A => n11690, ZN => n11694);
   U4980 : NAND2_X1 port map( A1 => n11692, A2 => n11691, ZN => n11693);
   U4981 : XNOR2_X1 port map( A => n11693, B => n11694, ZN => n11794);
   U4982 : MUX2_X1 port map( A => n13979, B => n13908, S => n11703, Z => n11697
                           );
   U4983 : MUX2_X1 port map( A => n14728, B => n13920, S => n10905, Z => n11695
                           );
   U4984 : INV_X1 port map( A => n11695, ZN => n11696);
   U4985 : NOR2_X1 port map( A1 => n11697, A2 => n11696, ZN => n11714);
   U4986 : MUX2_X1 port map( A => n11043, B => n10680, S => n8401, Z => n11699)
                           ;
   U4987 : MUX2_X1 port map( A => n10725, B => n11149, S => n10635, Z => n11698
                           );
   U4988 : NAND2_X1 port map( A1 => n11699, A2 => n11698, ZN => n11729);
   U4989 : MUX2_X1 port map( A => n14020, B => n10940, S => n11965, Z => n11701
                           );
   U4990 : NAND2_X1 port map( A1 => n14464, A2 => n12230, ZN => n11700);
   U4991 : NAND2_X1 port map( A1 => n11701, A2 => n11700, ZN => n11730);
   U4992 : NAND2_X1 port map( A1 => n11729, A2 => n11730, ZN => n11728);
   U4993 : NAND2_X1 port map( A1 => n11714, A2 => n11728, ZN => n12865);
   U4994 : INV_X1 port map( A => n12865, ZN => n11717);
   U4995 : XNOR2_X1 port map( A => n13368, B => n10873, ZN => n11702);
   U4996 : NAND2_X1 port map( A1 => n11702, A2 => n10679, ZN => n11706);
   U4997 : NAND2_X1 port map( A1 => n11704, A2 => n14737, ZN => n11705);
   U4998 : NAND2_X1 port map( A1 => n11706, A2 => n11705, ZN => n11712);
   U4999 : OAI21_X1 port map( B1 => n10977, B2 => n11707, A => n14833, ZN => 
                           n11711);
   U5000 : OR2_X1 port map( A1 => n11712, A2 => n11711, ZN => n12877);
   U5001 : MUX2_X1 port map( A => n10640, B => n13868, S => n14025, Z => n11710
                           );
   U5002 : XNOR2_X1 port map( A => n13265, B => n14593, ZN => n11708);
   U5003 : NAND2_X1 port map( A1 => n14813, A2 => n11708, ZN => n11709);
   U5004 : NAND2_X1 port map( A1 => n11710, A2 => n11709, ZN => n12878);
   U5005 : NAND2_X1 port map( A1 => n12877, A2 => n12878, ZN => n11713);
   U5006 : NAND2_X1 port map( A1 => n11712, A2 => n11711, ZN => n12876);
   U5007 : AND2_X1 port map( A1 => n11713, A2 => n12876, ZN => n12866);
   U5008 : INV_X1 port map( A => n11714, ZN => n11716);
   U5009 : INV_X1 port map( A => n11728, ZN => n11715);
   U5010 : NAND2_X1 port map( A1 => n11716, A2 => n11715, ZN => n12864);
   U5011 : XNOR2_X1 port map( A => n11719, B => n10741, ZN => n11720);
   U5012 : XNOR2_X1 port map( A => n11721, B => n11720, ZN => n11795);
   U5013 : XNOR2_X1 port map( A => n11795, B => n11792, ZN => n11722);
   U5014 : XNOR2_X1 port map( A => n11722, B => n11794, ZN => n13171);
   U5015 : MUX2_X1 port map( A => n13979, B => n12837, S => n13485, Z => n11725
                           );
   U5016 : MUX2_X1 port map( A => n13920, B => n14728, S => n14788, Z => n11723
                           );
   U5017 : INV_X1 port map( A => n11723, ZN => n11724);
   U5018 : NOR2_X1 port map( A1 => n11725, A2 => n11724, ZN => n11731);
   U5019 : MUX2_X1 port map( A => n13448, B => n13449, S => n14594, Z => n11727
                           );
   U5020 : MUX2_X1 port map( A => n14833, B => n13451, S => n14719, Z => n11726
                           );
   U5021 : AND2_X1 port map( A1 => n11727, A2 => n11726, ZN => n11732);
   U5022 : NAND2_X1 port map( A1 => n11731, A2 => n11732, ZN => n13180);
   U5023 : INV_X1 port map( A => n11731, ZN => n11734);
   U5024 : INV_X1 port map( A => n11732, ZN => n11733);
   U5025 : NAND2_X1 port map( A1 => n11734, A2 => n11733, ZN => n13179);
   U5026 : NAND2_X1 port map( A1 => n11735, A2 => n13179, ZN => n13174);
   U5027 : MUX2_X1 port map( A => n13448, B => n13449, S => n14025, Z => n11737
                           );
   U5028 : MUX2_X1 port map( A => n14833, B => n12783, S => n14777, Z => n11736
                           );
   U5029 : MUX2_X1 port map( A => n14017, B => n11201, S => n8351, Z => n11740)
                           ;
   U5030 : MUX2_X1 port map( A => n13915, B => n14779, S => n11738, Z => n11739
                           );
   U5031 : INV_X1 port map( A => n11761, ZN => n11741);
   U5032 : XNOR2_X1 port map( A => n11742, B => n11741, ZN => n11748);
   U5033 : MUX2_X1 port map( A => n11743, B => n13323, S => n13914, Z => n11746
                           );
   U5034 : MUX2_X1 port map( A => n10640, B => n13868, S => n14593, Z => n11744
                           );
   U5035 : INV_X1 port map( A => n11744, ZN => n11745);
   U5036 : NOR2_X1 port map( A1 => n11746, A2 => n11745, ZN => n11762);
   U5037 : INV_X1 port map( A => n11762, ZN => n11747);
   U5038 : XNOR2_X1 port map( A => n11748, B => n11747, ZN => n13173);
   U5039 : INV_X1 port map( A => n13173, ZN => n11756);
   U5040 : MUX2_X1 port map( A => n11043, B => n10680, S => n13924, Z => n11750
                           );
   U5041 : MUX2_X1 port map( A => n10725, B => n11834, S => n8401, Z => n11749)
                           ;
   U5042 : AND2_X1 port map( A1 => n11750, A2 => n11749, ZN => n11769);
   U5043 : INV_X1 port map( A => n11769, ZN => n11755);
   U5044 : AND2_X1 port map( A1 => n12174, A2 => n14719, ZN => n11765);
   U5045 : INV_X1 port map( A => n11765, ZN => n11753);
   U5046 : MUX2_X1 port map( A => n14020, B => n10939, S => n10914, Z => n11752
                           );
   U5047 : NAND2_X1 port map( A1 => n14457, A2 => n12230, ZN => n11751);
   U5048 : NAND2_X1 port map( A1 => n11752, A2 => n11751, ZN => n11766);
   U5049 : XNOR2_X1 port map( A => n11753, B => n11766, ZN => n11754);
   U5050 : XNOR2_X1 port map( A => n11755, B => n11754, ZN => n12862);
   U5051 : NAND2_X1 port map( A1 => n11756, A2 => n12862, ZN => n11757);
   U5052 : NAND2_X1 port map( A1 => n13174, A2 => n11757, ZN => n11759);
   U5053 : INV_X1 port map( A => n12862, ZN => n13172);
   U5054 : NAND2_X1 port map( A1 => n13173, A2 => n13172, ZN => n11758);
   U5055 : NAND2_X1 port map( A1 => n11759, A2 => n11758, ZN => n11778);
   U5056 : OAI21_X1 port map( B1 => n11762, B2 => n11761, A => n11760, ZN => 
                           n11764);
   U5057 : NAND2_X1 port map( A1 => n11762, A2 => n11761, ZN => n11763);
   U5058 : NAND2_X1 port map( A1 => n11764, A2 => n11763, ZN => n11782);
   U5059 : INV_X1 port map( A => n11782, ZN => n11777);
   U5060 : NAND2_X1 port map( A1 => n11766, A2 => n11765, ZN => n11768);
   U5061 : NOR2_X1 port map( A1 => n11766, A2 => n11765, ZN => n11767);
   U5062 : AOI21_X1 port map( B1 => n11769, B2 => n11768, A => n11767, ZN => 
                           n11773);
   U5063 : OAI21_X1 port map( B1 => n11771, B2 => n11770, A => n11786, ZN => 
                           n11774);
   U5064 : INV_X1 port map( A => n11774, ZN => n11772);
   U5065 : NAND2_X1 port map( A1 => n11773, A2 => n11772, ZN => n11781);
   U5066 : INV_X1 port map( A => n11773, ZN => n11775);
   U5067 : NAND2_X1 port map( A1 => n11775, A2 => n11774, ZN => n11783);
   U5068 : NAND2_X1 port map( A1 => n11781, A2 => n11783, ZN => n11776);
   U5069 : XNOR2_X1 port map( A => n11777, B => n11776, ZN => n13175);
   U5070 : OAI21_X1 port map( B1 => n13171, B2 => n11778, A => n13175, ZN => 
                           n11780);
   U5071 : NAND2_X1 port map( A1 => n13171, A2 => n11778, ZN => n11779);
   U5072 : NAND2_X1 port map( A1 => n11782, A2 => n11781, ZN => n11784);
   U5073 : NAND2_X1 port map( A1 => n11784, A2 => n11783, ZN => n11823);
   U5074 : XNOR2_X1 port map( A => n11790, B => n11820, ZN => n11791);
   U5075 : XNOR2_X1 port map( A => n11823, B => n11791, ZN => n11805);
   U5076 : NAND2_X1 port map( A1 => n11794, A2 => n11795, ZN => n11793);
   U5077 : NAND2_X1 port map( A1 => n11793, A2 => n11792, ZN => n11799);
   U5078 : INV_X1 port map( A => n11794, ZN => n11797);
   U5079 : INV_X1 port map( A => n11795, ZN => n11796);
   U5080 : NAND2_X1 port map( A1 => n11797, A2 => n11796, ZN => n11798);
   U5081 : NAND2_X1 port map( A1 => n11799, A2 => n11798, ZN => n11806);
   U5082 : INV_X1 port map( A => n11802, ZN => n11803);
   U5083 : XNOR2_X1 port map( A => n11806, B => n11804, ZN => n13525);
   U5084 : XOR2_X1 port map( A => n13525, B => n10906, Z => n11810);
   U5085 : OAI21_X1 port map( B1 => n11804, B2 => n11806, A => n11805, ZN => 
                           n11808);
   U5086 : NAND2_X1 port map( A1 => n11806, A2 => n11804, ZN => n11807);
   U5087 : INV_X1 port map( A => n13616, ZN => n11809);
   U5088 : NAND2_X1 port map( A1 => n11810, A2 => n11809, ZN => n11827);
   U5089 : NAND2_X1 port map( A1 => n11812, A2 => n11811, ZN => n11815);
   U5090 : INV_X1 port map( A => n11813, ZN => n11814);
   U5091 : XNOR2_X1 port map( A => n11815, B => n11814, ZN => n13896);
   U5092 : INV_X1 port map( A => n13896, ZN => n11818);
   U5093 : NAND2_X1 port map( A1 => n11817, A2 => n11816, ZN => n13893);
   U5094 : XNOR2_X1 port map( A => n11818, B => n13893, ZN => n11826);
   U5095 : NAND2_X1 port map( A1 => n11819, A2 => n11820, ZN => n11822);
   U5096 : NOR2_X1 port map( A1 => n11819, A2 => n11820, ZN => n11821);
   U5097 : AOI21_X1 port map( B1 => n11823, B2 => n11822, A => n11821, ZN => 
                           n13895);
   U5098 : INV_X1 port map( A => n13895, ZN => n11824);
   U5099 : XNOR2_X1 port map( A => n11824, B => n13891, ZN => n11825);
   U5100 : XNOR2_X1 port map( A => n11826, B => n11825, ZN => n13603);
   U5101 : OAI21_X1 port map( B1 => n10755, B2 => n10845, A => n10757, ZN => 
                           n14750);
   U5102 : INV_X1 port map( A => n11828, ZN => n11833);
   U5103 : NAND2_X1 port map( A1 => n11830, A2 => n11829, ZN => n11831);
   U5104 : MUX2_X1 port map( A => n14818, B => n11149, S => n12125, Z => n11835
                           );
   U5105 : MUX2_X1 port map( A => n10925, B => n10737, S => n14788, Z => n11839
                           );
   U5106 : XNOR2_X1 port map( A => n10905, B => n10693, ZN => n11837);
   U5107 : NAND2_X1 port map( A1 => n10971, A2 => n11837, ZN => n11838);
   U5110 : MUX2_X1 port map( A => n14878, B => n11971, S => n14465, Z => n11842
                           );
   U5111 : XNOR2_X1 port map( A => n14731, B => n10879, ZN => n11840);
   U5112 : NAND2_X1 port map( A1 => n14789, A2 => n11840, ZN => n11841);
   U5113 : NAND2_X1 port map( A1 => n11843, A2 => n12032, ZN => n11846);
   U5114 : MUX2_X1 port map( A => n13817, B => n10885, S => n13914, Z => n11845
                           );
   U5115 : MUX2_X1 port map( A => n11995, B => n14882, S => n14785, Z => n11844
                           );
   U5116 : NAND2_X1 port map( A1 => n11845, A2 => n11844, ZN => n11847);
   U5117 : OAI211_X1 port map( C1 => n12034, C2 => n12033, A => n11846, B => 
                           n11847, ZN => n13030);
   U5118 : INV_X1 port map( A => n12032, ZN => n11848);
   U5119 : OAI21_X1 port map( B1 => n12034, B2 => n11848, A => n12033, ZN => 
                           n11850);
   U5120 : AOI21_X1 port map( B1 => n12034, B2 => n11848, A => n11847, ZN => 
                           n11849);
   U5121 : NAND2_X1 port map( A1 => n13030, A2 => n13028, ZN => n11856);
   U5122 : MUX2_X1 port map( A => n13283, B => n14716, S => n10914, Z => n11912
                           );
   U5123 : NOR2_X1 port map( A1 => n14594, A2 => n13482, ZN => n11909);
   U5124 : NAND2_X1 port map( A1 => n11909, A2 => n14784, ZN => n11851);
   U5125 : AND2_X1 port map( A1 => n11912, A2 => n11851, ZN => n11852);
   U5126 : MUX2_X1 port map( A => n13346, B => n12805, S => n10743, Z => n11913
                           );
   U5127 : NAND2_X1 port map( A1 => n11852, A2 => n11913, ZN => n11855);
   U5128 : INV_X1 port map( A => n11909, ZN => n11853);
   U5129 : NAND2_X1 port map( A1 => n11853, A2 => n11594, ZN => n11854);
   U5130 : NAND2_X1 port map( A1 => n11855, A2 => n11854, ZN => n13026);
   U5131 : XNOR2_X1 port map( A => n11856, B => n13026, ZN => n14084);
   U5132 : MUX2_X1 port map( A => n13442, B => n10737, S => n14448, Z => n11858
                           );
   U5133 : NAND2_X1 port map( A1 => n11857, A2 => n13279, ZN => n11860);
   U5134 : NAND2_X1 port map( A1 => n11858, A2 => n11860, ZN => n11954);
   U5135 : NOR2_X1 port map( A1 => n10864, A2 => n13482, ZN => n11951);
   U5136 : NAND2_X1 port map( A1 => n11954, A2 => n11951, ZN => n11868);
   U5137 : INV_X1 port map( A => n11858, ZN => n11866);
   U5138 : INV_X1 port map( A => n11951, ZN => n11859);
   U5139 : NAND2_X1 port map( A1 => n11860, A2 => n11859, ZN => n11865);
   U5140 : MUX2_X1 port map( A => n13347, B => n14716, S => n12743, Z => n11864
                           );
   U5141 : XNOR2_X1 port map( A => n10913, B => n11861, ZN => n11862);
   U5142 : NAND2_X1 port map( A1 => n12174, A2 => n11862, ZN => n11863);
   U5143 : NAND2_X1 port map( A1 => n11864, A2 => n11863, ZN => n11952);
   U5144 : OAI21_X1 port map( B1 => n11866, B2 => n11865, A => n11952, ZN => 
                           n11867);
   U5145 : NAND2_X1 port map( A1 => n11867, A2 => n11868, ZN => n11921);
   U5146 : MUX2_X1 port map( A => n10885, B => n14880, S => n14593, Z => n11870
                           );
   U5147 : MUX2_X1 port map( A => n13819, B => n14882, S => n14447, Z => n11869
                           );
   U5148 : NAND2_X1 port map( A1 => n11870, A2 => n11869, ZN => n11920);
   U5149 : NAND2_X1 port map( A1 => n11921, A2 => n11920, ZN => n11878);
   U5150 : MUX2_X1 port map( A => n14878, B => n11971, S => n14593, Z => n11871
                           );
   U5151 : NAND2_X1 port map( A1 => n11872, A2 => n11871, ZN => n11993);
   U5152 : AOI21_X1 port map( B1 => n14501, B2 => n14881, A => n14586, ZN => 
                           n11922);
   U5153 : MUX2_X1 port map( A => n10725, B => n11834, S => n13810, Z => n11875
                           );
   U5154 : XOR2_X1 port map( A => n8329, B => n14717, Z => n11873);
   U5155 : NAND2_X1 port map( A1 => n11873, A2 => n10857, ZN => n11874);
   U5156 : NAND2_X1 port map( A1 => n11875, A2 => n11874, ZN => n11992);
   U5157 : OAI21_X1 port map( B1 => n11993, B2 => n11922, A => n11992, ZN => 
                           n11877);
   U5158 : NAND2_X1 port map( A1 => n11993, A2 => n11922, ZN => n11876);
   U5159 : NAND3_X1 port map( A1 => n11878, A2 => n11877, A3 => n11876, ZN => 
                           n11882);
   U5160 : INV_X1 port map( A => n11921, ZN => n11880);
   U5161 : INV_X1 port map( A => n11920, ZN => n11879);
   U5162 : NAND2_X1 port map( A1 => n11880, A2 => n11879, ZN => n11881);
   U5163 : NAND2_X1 port map( A1 => n11882, A2 => n11881, ZN => n14083);
   U5164 : MUX2_X1 port map( A => n11096, B => n12837, S => n13450, Z => n11885
                           );
   U5165 : MUX2_X1 port map( A => n13980, B => n14728, S => n10726, Z => n11883
                           );
   U5166 : INV_X1 port map( A => n11883, ZN => n11884);
   U5167 : OR2_X2 port map( A1 => n11885, A2 => n11884, ZN => n11988);
   U5168 : MUX2_X1 port map( A => n14833, B => n12783, S => n10743, Z => n11888
                           );
   U5169 : XNOR2_X1 port map( A => n14725, B => n10869, ZN => n11886);
   U5170 : NAND2_X1 port map( A1 => n14727, A2 => n11886, ZN => n11887);
   U5171 : NAND2_X1 port map( A1 => n11888, A2 => n11887, ZN => n11987);
   U5172 : NAND2_X1 port map( A1 => n11988, A2 => n11987, ZN => n11891);
   U5173 : MUX2_X1 port map( A => n13323, B => n11743, S => n10831, Z => n11890
                           );
   U5174 : MUX2_X1 port map( A => n11385, B => n11933, S => n14452, Z => n11889
                           );
   U5175 : NAND2_X1 port map( A1 => n11891, A2 => n11989, ZN => n11895);
   U5176 : INV_X1 port map( A => n11988, ZN => n11893);
   U5177 : INV_X1 port map( A => n11987, ZN => n11892);
   U5178 : NAND2_X1 port map( A1 => n11893, A2 => n11892, ZN => n11894);
   U5179 : NAND2_X1 port map( A1 => n11895, A2 => n11894, ZN => n14088);
   U5180 : MUX2_X1 port map( A => n14114, B => n13362, S => B_SIG_8_port, Z => 
                           n11899);
   U5181 : NAND2_X1 port map( A1 => n11225, A2 => n10904, ZN => n11897);
   U5182 : NAND2_X1 port map( A1 => n12146, A2 => n14451, ZN => n11896);
   U5183 : NAND2_X1 port map( A1 => n11897, A2 => n11896, ZN => n11898);
   U5185 : MUX2_X1 port map( A => n13373, B => n10641, S => n13368, Z => n12916
                           );
   U5186 : MUX2_X1 port map( A => n13372, B => n13371, S => n8351, Z => n12917)
                           ;
   U5187 : NAND3_X1 port map( A1 => n12915, A2 => n12916, A3 => n12917, ZN => 
                           n11904);
   U5188 : MUX2_X1 port map( A => n11900, B => n11201, S => n14117, Z => n11902
                           );
   U5189 : MUX2_X1 port map( A => n13915, B => n14779, S => n8334, Z => n11901)
                           ;
   U5190 : NAND2_X1 port map( A1 => n11902, A2 => n11901, ZN => n12914);
   U5191 : NAND2_X1 port map( A1 => n12915, A2 => n11905, ZN => n11903);
   U5192 : AND2_X1 port map( A1 => n11903, A2 => n11904, ZN => n11908);
   U5193 : INV_X1 port map( A => n12914, ZN => n11905);
   U5194 : AND2_X1 port map( A1 => n11905, A2 => n12916, ZN => n11906);
   U5195 : NAND2_X1 port map( A1 => n12917, A2 => n11906, ZN => n11907);
   U5196 : XNOR2_X1 port map( A => n11909, B => n11594, ZN => n11911);
   U5197 : AOI21_X1 port map( B1 => n11913, B2 => n11912, A => n11911, ZN => 
                           n11910);
   U5198 : INV_X1 port map( A => n11910, ZN => n11915);
   U5199 : NAND3_X1 port map( A1 => n11913, A2 => n11912, A3 => n11911, ZN => 
                           n11914);
   U5200 : NAND2_X1 port map( A1 => n11915, A2 => n11914, ZN => n11916);
   U5201 : NAND2_X1 port map( A1 => n12007, A2 => n11916, ZN => n14087);
   U5202 : NAND2_X1 port map( A1 => n14088, A2 => n14087, ZN => n11918);
   U5203 : INV_X1 port map( A => n11916, ZN => n12008);
   U5204 : INV_X1 port map( A => n12007, ZN => n11917);
   U5205 : NAND2_X1 port map( A1 => n12008, A2 => n11917, ZN => n14086);
   U5206 : NAND2_X1 port map( A1 => n11918, A2 => n14086, ZN => n14085);
   U5207 : XNOR2_X1 port map( A => n11921, B => n11920, ZN => n11927);
   U5208 : INV_X1 port map( A => n11993, ZN => n11925);
   U5209 : NAND2_X1 port map( A1 => n11992, A2 => n11922, ZN => n11924);
   U5210 : INV_X1 port map( A => n11992, ZN => n11923);
   U5211 : INV_X1 port map( A => n11922, ZN => n11991);
   U5212 : AOI22_X1 port map( A1 => n11925, A2 => n11924, B1 => n11923, B2 => 
                           n11991, ZN => n11926);
   U5213 : XNOR2_X1 port map( A => n11927, B => n11926, ZN => n13133);
   U5214 : INV_X1 port map( A => n14466, ZN => n13282);
   U5215 : MUX2_X1 port map( A => n11096, B => n13908, S => n13282, Z => n11930
                           );
   U5216 : MUX2_X1 port map( A => n13920, B => n14728, S => n14450, Z => n11928
                           );
   U5217 : INV_X1 port map( A => n11928, ZN => n11929);
   U5218 : NOR2_X1 port map( A1 => n11930, A2 => n11929, ZN => n13067);
   U5219 : MUX2_X1 port map( A => n11743, B => n13323, S => n13234, Z => n11938
                           );
   U5220 : MUX2_X1 port map( A => n13372, B => n13371, S => n13368, Z => n11932
                           );
   U5221 : MUX2_X1 port map( A => n10745, B => n13373, S => n14819, Z => n11931
                           );
   U5222 : NAND2_X1 port map( A1 => n11932, A2 => n11931, ZN => n11939);
   U5223 : NAND2_X1 port map( A1 => n11938, A2 => n11939, ZN => n11936);
   U5224 : NAND2_X1 port map( A1 => n11939, A2 => n11937, ZN => n11935);
   U5225 : NAND3_X1 port map( A1 => n13067, A2 => n11936, A3 => n11935, ZN => 
                           n11941);
   U5226 : NOR2_X1 port map( A1 => n11938, A2 => n11937, ZN => n13069);
   U5227 : INV_X1 port map( A => n11939, ZN => n13068);
   U5228 : NAND2_X1 port map( A1 => n13069, A2 => n13068, ZN => n11940);
   U5229 : NAND2_X1 port map( A1 => n11941, A2 => n11940, ZN => n13084);
   U5230 : INV_X1 port map( A => n14467, ZN => n13262);
   U5231 : MUX2_X1 port map( A => n14017, B => n11201, S => n13262, Z => n11943
                           );
   U5232 : MUX2_X1 port map( A => n13915, B => n14779, S => n13450, Z => n11942
                           );
   U5233 : NAND2_X1 port map( A1 => n11943, A2 => n11942, ZN => n13106);
   U5234 : NAND2_X1 port map( A1 => n10630, A2 => n10904, ZN => n11944);
   U5235 : OAI21_X1 port map( B1 => n14114, B2 => n10904, A => n11944, ZN => 
                           n11946);
   U5236 : MUX2_X1 port map( A => n10713, B => n10636, S => n13924, Z => n11945
                           );
   U5237 : NAND2_X1 port map( A1 => n11946, A2 => n11945, ZN => n13107);
   U5238 : MUX2_X1 port map( A => n13449, B => n13448, S => n10743, Z => n11948
                           );
   U5239 : MUX2_X1 port map( A => n14833, B => n12783, S => n10914, Z => n11947
                           );
   U5240 : NAND2_X1 port map( A1 => n11948, A2 => n11947, ZN => n13115);
   U5241 : OAI21_X1 port map( B1 => n13106, B2 => n13107, A => n13115, ZN => 
                           n11950);
   U5242 : NAND2_X1 port map( A1 => n13106, A2 => n13107, ZN => n11949);
   U5243 : AND2_X1 port map( A1 => n11950, A2 => n11949, ZN => n13085);
   U5244 : OR2_X1 port map( A1 => n13084, A2 => n13085, ZN => n11956);
   U5245 : XNOR2_X1 port map( A => n10730, B => n11951, ZN => n11953);
   U5246 : XOR2_X1 port map( A => n11954, B => n11953, Z => n13086);
   U5247 : AND2_X1 port map( A1 => n13084, A2 => n13085, ZN => n11955);
   U5248 : NOR2_X1 port map( A1 => n13133, A2 => n13134, ZN => n11986);
   U5249 : MUX2_X1 port map( A => n11043, B => n10680, S => n13810, Z => n11959
                           );
   U5250 : MUX2_X1 port map( A => n10725, B => n11149, S => n14478, Z => n11958
                           );
   U5251 : NAND2_X1 port map( A1 => n11959, A2 => n11958, ZN => n13109);
   U5252 : MUX2_X1 port map( A => n10925, B => n10738, S => n14465, Z => n11962
                           );
   U5253 : XOR2_X1 port map( A => n13277, B => n8401, Z => n11960);
   U5254 : NAND2_X1 port map( A1 => n10971, A2 => n11960, ZN => n11961);
   U5255 : NAND2_X1 port map( A1 => n11962, A2 => n11961, ZN => n13111);
   U5256 : MUX2_X1 port map( A => n10885, B => n14880, S => n14025, Z => n11964
                           );
   U5257 : MUX2_X1 port map( A => n13819, B => n14882, S => n14777, Z => n11963
                           );
   U5258 : NAND2_X1 port map( A1 => n11964, A2 => n11963, ZN => n11981);
   U5259 : NAND2_X1 port map( A1 => n12922, A2 => n11981, ZN => n11980);
   U5260 : MUX2_X1 port map( A => n13283, B => n14716, S => n8351, Z => n11968)
                           ;
   U5261 : XNOR2_X1 port map( A => n11965, B => n10877, ZN => n11966);
   U5262 : NAND2_X1 port map( A1 => n11966, A2 => n12174, ZN => n11967);
   U5263 : NAND2_X1 port map( A1 => n11968, A2 => n11967, ZN => n11975);
   U5264 : MUX2_X1 port map( A => n10939, B => n14020, S => n10841, Z => n11970
                           );
   U5265 : NAND2_X1 port map( A1 => n14459, A2 => n12230, ZN => n11969);
   U5266 : NAND2_X1 port map( A1 => n11970, A2 => n11969, ZN => n11976);
   U5267 : NAND2_X1 port map( A1 => n11975, A2 => n11976, ZN => n13076);
   U5268 : MUX2_X1 port map( A => n13824, B => n11971, S => n14025, Z => n11974
                           );
   U5269 : XNOR2_X1 port map( A => n14785, B => n10879, ZN => n11972);
   U5270 : NAND2_X1 port map( A1 => n14789, A2 => n11972, ZN => n11973);
   U5271 : AND2_X1 port map( A1 => n11974, A2 => n11973, ZN => n13078);
   U5272 : NAND2_X1 port map( A1 => n13076, A2 => n13078, ZN => n11979);
   U5273 : INV_X1 port map( A => n11975, ZN => n11978);
   U5274 : INV_X1 port map( A => n11976, ZN => n11977);
   U5275 : NAND2_X1 port map( A1 => n11978, A2 => n11977, ZN => n13077);
   U5276 : NAND2_X1 port map( A1 => n11979, A2 => n13077, ZN => n12923);
   U5277 : NAND2_X1 port map( A1 => n11980, A2 => n12923, ZN => n11984);
   U5278 : INV_X1 port map( A => n12922, ZN => n11982);
   U5279 : INV_X1 port map( A => n11981, ZN => n12921);
   U5280 : NAND2_X1 port map( A1 => n11982, A2 => n12921, ZN => n11983);
   U5281 : NAND2_X1 port map( A1 => n11984, A2 => n11983, ZN => n13132);
   U5282 : NAND2_X1 port map( A1 => n13134, A2 => n13133, ZN => n11985);
   U5283 : OAI21_X2 port map( B1 => n11986, B2 => n13132, A => n11985, ZN => 
                           n13551);
   U5284 : XNOR2_X1 port map( A => n13221, B => n13551, ZN => n14809);
   U5285 : XNOR2_X1 port map( A => n11988, B => n11987, ZN => n11990);
   U5286 : XNOR2_X1 port map( A => n11990, B => n11989, ZN => n12004);
   U5287 : XNOR2_X1 port map( A => n11992, B => n11991, ZN => n11994);
   U5288 : XNOR2_X1 port map( A => n11994, B => n11993, ZN => n12005);
   U5289 : NAND2_X1 port map( A1 => n12004, A2 => n12005, ZN => n12927);
   U5290 : XNOR2_X1 port map( A => n13109, B => n10915, ZN => n11999);
   U5291 : INV_X1 port map( A => n11995, ZN => n13486);
   U5292 : AOI21_X1 port map( B1 => n14487, B2 => n10864, A => n13486, ZN => 
                           n13110);
   U5293 : NAND2_X1 port map( A1 => n11999, A2 => n13110, ZN => n11998);
   U5294 : MUX2_X1 port map( A => n10885, B => n13817, S => n14594, Z => n11997
                           );
   U5295 : MUX2_X1 port map( A => n13819, B => n14882, S => n14719, Z => n11996
                           );
   U5296 : NAND2_X1 port map( A1 => n11997, A2 => n11996, ZN => n13108);
   U5297 : NAND2_X1 port map( A1 => n11998, A2 => n13108, ZN => n12003);
   U5298 : INV_X1 port map( A => n11999, ZN => n12001);
   U5299 : INV_X1 port map( A => n13110, ZN => n12000);
   U5300 : NAND2_X1 port map( A1 => n12001, A2 => n12000, ZN => n12002);
   U5301 : NAND2_X1 port map( A1 => n12003, A2 => n12002, ZN => n12928);
   U5302 : NAND2_X1 port map( A1 => n12927, A2 => n12928, ZN => n12006);
   U5303 : NAND2_X1 port map( A1 => n12006, A2 => n12926, ZN => n13187);
   U5304 : XNOR2_X1 port map( A => n14088, B => n12007, ZN => n12009);
   U5305 : XNOR2_X1 port map( A => n12009, B => n12008, ZN => n13189);
   U5306 : MUX2_X1 port map( A => n10640, B => n13868, S => n10831, Z => n12013
                           );
   U5307 : XNOR2_X1 port map( A => n12010, B => n13813, ZN => n12011);
   U5308 : NAND2_X1 port map( A1 => n14813, A2 => n12011, ZN => n12012);
   U5309 : MUX2_X1 port map( A => n14728, B => n13980, S => n13450, Z => n12017
                           );
   U5310 : XNOR2_X1 port map( A => n12014, B => n8334, ZN => n12015);
   U5311 : NAND2_X1 port map( A1 => n14786, A2 => n12015, ZN => n12016);
   U5312 : NAND2_X1 port map( A1 => n12017, A2 => n12016, ZN => n13017);
   U5313 : XNOR2_X1 port map( A => n13017, B => n13013, ZN => n12022);
   U5314 : MUX2_X1 port map( A => n14833, B => n12783, S => n14449, Z => n12021
                           );
   U5315 : XNOR2_X1 port map( A => n12018, B => n12246, ZN => n12019);
   U5316 : NAND2_X1 port map( A1 => n12019, A2 => n14727, ZN => n12020);
   U5317 : NAND2_X1 port map( A1 => n12021, A2 => n12020, ZN => n13016);
   U5318 : XNOR2_X1 port map( A => n12022, B => n13016, ZN => n13140);
   U5319 : INV_X1 port map( A => n13140, ZN => n13143);
   U5320 : MUX2_X1 port map( A => n14456, B => n14779, S => n14117, Z => n12025
                           );
   U5321 : XNOR2_X1 port map( A => FP_A(3), B => n14646, ZN => n10840);
   U5322 : NAND2_X1 port map( A1 => n10679, A2 => n12023, ZN => n12024);
   U5323 : NAND2_X1 port map( A1 => n12025, A2 => n12024, ZN => n13005);
   U5324 : MUX2_X1 port map( A => n12142, B => n10745, S => n8351, Z => n12027)
                           ;
   U5325 : XNOR2_X1 port map( A => n8392, B => n12671, ZN => n12026);
   U5326 : NAND2_X1 port map( A1 => n12026, A2 => n12640, ZN => n13002);
   U5327 : XNOR2_X1 port map( A => n13005, B => n13006, ZN => n12031);
   U5328 : MUX2_X1 port map( A => n14114, B => n13362, S => n13368, Z => n12029
                           );
   U5329 : MUX2_X1 port map( A => n12146, B => n11225, S => B_SIG_8_port, Z => 
                           n12028);
   U5330 : XNOR2_X1 port map( A => n12031, B => n12030, ZN => n13141);
   U5331 : XNOR2_X1 port map( A => n12033, B => n12032, ZN => n12035);
   U5332 : XNOR2_X1 port map( A => n13141, B => n13144, ZN => n12036);
   U5333 : XNOR2_X1 port map( A => n12036, B => n13143, ZN => n13188);
   U5334 : OAI21_X1 port map( B1 => n13187, B2 => n13189, A => n13188, ZN => 
                           n12041);
   U5335 : INV_X1 port map( A => n12928, ZN => n12037);
   U5336 : NAND2_X1 port map( A1 => n12926, A2 => n12037, ZN => n12038);
   U5337 : NAND3_X1 port map( A1 => n13189, A2 => n12927, A3 => n12038, ZN => 
                           n12040);
   U5338 : NAND2_X1 port map( A1 => n12040, A2 => n12041, ZN => n14811);
   U5339 : XNOR2_X1 port map( A => n14809, B => n10727, ZN => n14792);
   U5340 : INV_X1 port map( A => FP_B(6), ZN => n14557);
   U5341 : INV_X1 port map( A => FP_A(17), ZN => n14671);
   U5342 : INV_X1 port map( A => FP_A(11), ZN => n14698);
   U5344 : INV_X1 port map( A => FP_A(15), ZN => n384);
   U5345 : AND2_X1 port map( A1 => FP_A(11), A2 => n14667, ZN => n14668);
   U5346 : AND2_X1 port map( A1 => FP_A(17), A2 => FP_A(18), ZN => n14709);
   U5347 : INV_X1 port map( A => n14709, ZN => n14639);
   U5348 : INV_X1 port map( A => FP_A(8), ZN => n14708);
   U5349 : INV_X1 port map( A => FP_B(8), ZN => n14591);
   U5350 : INV_X1 port map( A => FP_A(4), ZN => n14702);
   U5351 : NOR2_X1 port map( A1 => FP_A(6), A2 => FP_A(5), ZN => n12068);
   U5352 : INV_X1 port map( A => n12068, ZN => n14524);
   U5353 : INV_X1 port map( A => FP_A(2), ZN => n12047);
   U5354 : OR2_X1 port map( A1 => n12047, A2 => n12567, ZN => n12048);
   U5355 : OR2_X1 port map( A1 => FP_A(3), A2 => n12048, ZN => n14672);
   U5356 : NOR2_X1 port map( A1 => FP_A(22), A2 => FP_A(21), ZN => n12064);
   U5357 : INV_X1 port map( A => n12064, ZN => n14523);
   U5358 : NAND2_X1 port map( A1 => FP_A(21), A2 => FP_A(22), ZN => n14663);
   U5359 : MUX2_X1 port map( A => n2593, B => n2592, S => n14729, Z => n14900);
   U5360 : INV_X1 port map( A => n14900, ZN => n14899);
   U5361 : MUX2_X1 port map( A => n2589, B => n8375, S => SIG_in_27_port, Z => 
                           n12049);
   U5362 : INV_X1 port map( A => n12049, ZN => n14918);
   U5363 : MUX2_X1 port map( A => n14521, B => n2590, S => SIG_in_27_port, Z =>
                           n14909);
   U5364 : INV_X1 port map( A => n14909, ZN => n14902);
   U5365 : NOR2_X1 port map( A1 => FP_B(24), A2 => FP_B(23), ZN => n12053);
   U5366 : NOR2_X1 port map( A1 => FP_B(26), A2 => FP_B(25), ZN => n12052);
   U5367 : NOR2_X1 port map( A1 => FP_B(28), A2 => FP_B(27), ZN => n12051);
   U5368 : NOR2_X1 port map( A1 => FP_B(30), A2 => FP_B(29), ZN => n12050);
   U5369 : NAND4_X1 port map( A1 => n12053, A2 => n12052, A3 => n12051, A4 => 
                           n12050, ZN => I1_I1_N13);
   U5370 : NOR2_X1 port map( A1 => FP_A(18), A2 => FP_A(17), ZN => n14732);
   U5371 : NOR2_X1 port map( A1 => FP_A(8), A2 => FP_A(7), ZN => n14733);
   U5372 : NOR2_X1 port map( A1 => FP_A(24), A2 => FP_A(23), ZN => n12057);
   U5373 : NOR2_X1 port map( A1 => FP_A(26), A2 => FP_A(25), ZN => n12056);
   U5374 : NOR2_X1 port map( A1 => FP_A(28), A2 => FP_A(27), ZN => n12055);
   U5375 : NOR2_X1 port map( A1 => FP_A(30), A2 => FP_A(29), ZN => n12054);
   U5376 : NAND4_X1 port map( A1 => n12057, A2 => n12056, A3 => n12055, A4 => 
                           n12054, ZN => I1_I0_N13);
   U5377 : NOR2_X1 port map( A1 => FP_A(16), A2 => FP_A(15), ZN => n12061);
   U5378 : NOR2_X1 port map( A1 => FP_A(14), A2 => FP_A(13), ZN => n12060);
   U5379 : NOR2_X1 port map( A1 => FP_A(12), A2 => FP_A(11), ZN => n12059);
   U5380 : NOR2_X1 port map( A1 => FP_A(10), A2 => FP_A(9), ZN => n12058);
   U5381 : NAND4_X1 port map( A1 => n12061, A2 => n12060, A3 => n12059, A4 => 
                           n12058, ZN => n12066);
   U5382 : NOR2_X1 port map( A1 => FP_A(20), A2 => FP_A(19), ZN => n12063);
   U5383 : INV_X1 port map( A => FP_A(0), ZN => n12062);
   U5384 : NAND4_X1 port map( A1 => n12064, A2 => n12063, A3 => n14732, A4 => 
                           n12062, ZN => n12065);
   U5385 : NOR2_X1 port map( A1 => n12066, A2 => n12065, ZN => n12070);
   U5386 : NOR2_X1 port map( A1 => FP_A(4), A2 => FP_A(3), ZN => n12067);
   U5387 : NOR2_X1 port map( A1 => FP_A(2), A2 => FP_A(1), ZN => n12334);
   U5388 : AND4_X1 port map( A1 => n14733, A2 => n12068, A3 => n12067, A4 => 
                           n12334, ZN => n12069);
   U5389 : AND2_X1 port map( A1 => n12070, A2 => n12069, ZN => n13844);
   U5390 : NAND4_X1 port map( A1 => FP_A(24), A2 => FP_A(23), A3 => FP_A(26), 
                           A4 => FP_A(25), ZN => n12072);
   U5391 : NAND4_X1 port map( A1 => FP_A(28), A2 => FP_A(27), A3 => FP_A(30), 
                           A4 => FP_A(29), ZN => n12071);
   U5392 : NOR2_X1 port map( A1 => n12072, A2 => n12071, ZN => n14419);
   U5393 : NAND2_X1 port map( A1 => n13844, A2 => n14419, ZN => n14422);
   U5394 : NOR2_X1 port map( A1 => FP_B(8), A2 => FP_B(7), ZN => n12076);
   U5395 : NOR2_X1 port map( A1 => FP_B(6), A2 => FP_B(5), ZN => n12075);
   U5396 : NOR2_X1 port map( A1 => FP_B(4), A2 => FP_B(3), ZN => n12074);
   U5397 : NOR2_X1 port map( A1 => FP_B(2), A2 => FP_B(1), ZN => n12073);
   U5398 : AND4_X1 port map( A1 => n12076, A2 => n12075, A3 => n12074, A4 => 
                           n12073, ZN => n12086);
   U5399 : NOR2_X1 port map( A1 => FP_B(16), A2 => FP_B(15), ZN => n12080);
   U5400 : NOR2_X1 port map( A1 => FP_B(14), A2 => FP_B(13), ZN => n12079);
   U5401 : NOR2_X1 port map( A1 => FP_B(12), A2 => FP_B(11), ZN => n12078);
   U5402 : NOR2_X1 port map( A1 => FP_B(10), A2 => FP_B(9), ZN => n12077);
   U5403 : AND4_X1 port map( A1 => n12080, A2 => n12079, A3 => n12078, A4 => 
                           n12077, ZN => n12085);
   U5404 : NOR3_X1 port map( A1 => FP_B(0), A2 => FP_B(22), A3 => FP_B(21), ZN 
                           => n12084);
   U5405 : NOR2_X1 port map( A1 => FP_B(20), A2 => FP_B(19), ZN => n12082);
   U5406 : NOR2_X1 port map( A1 => FP_B(18), A2 => FP_B(17), ZN => n12081);
   U5407 : AND2_X1 port map( A1 => n12082, A2 => n12081, ZN => n12083);
   U5408 : NAND4_X1 port map( A1 => n12086, A2 => n12085, A3 => n12084, A4 => 
                           n12083, ZN => n14421);
   U5409 : INV_X1 port map( A => n14421, ZN => n12092);
   U5410 : NAND4_X1 port map( A1 => FP_B(24), A2 => FP_B(23), A3 => FP_B(26), 
                           A4 => FP_B(25), ZN => n12088);
   U5411 : NAND4_X1 port map( A1 => FP_B(28), A2 => FP_B(27), A3 => FP_B(30), 
                           A4 => FP_B(29), ZN => n12087);
   U5412 : NOR2_X1 port map( A1 => n12088, A2 => n12087, ZN => n14423);
   U5413 : NAND2_X1 port map( A1 => n12092, A2 => n14423, ZN => n12089);
   U5414 : NAND2_X1 port map( A1 => n14422, A2 => n12089, ZN => n12094);
   U5415 : INV_X1 port map( A => I1_I0_N13, ZN => n13843);
   U5416 : NAND2_X1 port map( A1 => n13843, A2 => n14423, ZN => n12091);
   U5417 : INV_X1 port map( A => n13844, ZN => n14420);
   U5418 : INV_X1 port map( A => n14419, ZN => n12090);
   U5419 : OAI22_X1 port map( A1 => n12091, A2 => n14420, B1 => n12090, B2 => 
                           I1_I1_N13, ZN => n12093);
   U5420 : NAND2_X1 port map( A1 => n12093, A2 => n12092, ZN => n14426);
   U5421 : AND2_X1 port map( A1 => n12094, A2 => n14426, ZN => I1_isINF_int);
   U5422 : OAI21_X1 port map( B1 => n12095, B2 => n10942, A => n14328, ZN => 
                           n12096);
   U5423 : INV_X1 port map( A => n12096, ZN => I3_SIG_out_7_port);
   U5424 : NAND2_X1 port map( A1 => n12098, A2 => n12097, ZN => n12099);
   U5425 : AND2_X1 port map( A1 => n14338, A2 => n12099, ZN => 
                           I3_SIG_out_12_port);
   U5426 : XNOR2_X1 port map( A => n12342, B => n14690, ZN => n14429);
   U5427 : INV_X1 port map( A => n14429, ZN => n14921);
   U5429 : OAI21_X1 port map( B1 => n12265, B2 => n10758, A => n10789, ZN => 
                           n12101);
   U5430 : MUX2_X1 port map( A => n12631, B => n12102, S => n14881, Z => n12212
                           );
   U5431 : AND2_X1 port map( A1 => n13450, A2 => n13809, ZN => n12210);
   U5432 : INV_X1 port map( A => n12210, ZN => n12116);
   U5433 : MUX2_X1 port map( A => n14880, B => n10886, S => n13261, Z => n12104
                           );
   U5435 : MUX2_X1 port map( A => n13819, B => n14882, S => n8334, Z => n12103)
                           ;
   U5436 : NAND2_X1 port map( A1 => n12104, A2 => n12103, ZN => n12211);
   U5437 : OAI21_X1 port map( B1 => n12212, B2 => n12116, A => n12211, ZN => 
                           n12106);
   U5438 : NAND2_X1 port map( A1 => n12212, A2 => n12116, ZN => n12105);
   U5439 : NAND2_X1 port map( A1 => n12106, A2 => n12105, ZN => n12226);
   U5440 : NAND2_X1 port map( A1 => n13262, A2 => n13809, ZN => n12115);
   U5441 : XNOR2_X1 port map( A => n12116, B => n12115, ZN => n12107);
   U5442 : XNOR2_X1 port map( A => n12631, B => n12107, ZN => n12224);
   U5443 : MUX2_X1 port map( A => n10886, B => n14880, S => n10841, Z => n12109
                           );
   U5444 : MUX2_X1 port map( A => n13819, B => n14882, S => n13261, Z => n12108
                           );
   U5445 : NAND2_X1 port map( A1 => n12109, A2 => n12108, ZN => n12223);
   U5446 : INV_X1 port map( A => n12223, ZN => n12110);
   U5447 : NAND2_X1 port map( A1 => n12224, A2 => n12110, ZN => n12111);
   U5448 : NAND2_X1 port map( A1 => n12226, A2 => n12111, ZN => n12114);
   U5449 : INV_X1 port map( A => n12224, ZN => n12112);
   U5450 : NAND2_X1 port map( A1 => n12112, A2 => n12223, ZN => n12113);
   U5451 : NAND2_X1 port map( A1 => n12114, A2 => n12113, ZN => n14306);
   U5452 : AOI21_X1 port map( B1 => n12631, B2 => n12116, A => n12115, ZN => 
                           n12118);
   U5453 : NOR2_X1 port map( A1 => n12631, A2 => n12116, ZN => n12117);
   U5454 : NOR2_X1 port map( A1 => n12118, A2 => n12117, ZN => n14307);
   U5455 : OAI21_X1 port map( B1 => n13819, B2 => n14881, A => n14880, ZN => 
                           n12121);
   U5456 : AND2_X1 port map( A1 => n13261, A2 => n10702, ZN => n12119);
   U5457 : NOR2_X1 port map( A1 => n12121, A2 => n12119, ZN => n14300);
   U5458 : OR2_X1 port map( A1 => n14882, A2 => n10841, ZN => n12120);
   U5459 : AND2_X1 port map( A1 => n14300, A2 => n12120, ZN => n14298);
   U5460 : INV_X1 port map( A => n14298, ZN => n12122);
   U5461 : NAND2_X1 port map( A1 => n12121, A2 => n8331, ZN => n14309);
   U5462 : NAND2_X1 port map( A1 => n12122, A2 => n14309, ZN => n12123);
   U5463 : XNOR2_X1 port map( A => n14307, B => n12123, ZN => n14305);
   U5464 : INV_X1 port map( A => n14305, ZN => n14302);
   U5465 : XNOR2_X1 port map( A => n14306, B => n14302, ZN => n14914);
   U5466 : XOR2_X1 port map( A => n12124, B => n12125, Z => n12126);
   U5467 : NAND2_X1 port map( A1 => n12126, A2 => n14813, ZN => n12131);
   U5468 : NAND2_X1 port map( A1 => n10640, A2 => n13810, ZN => n12129);
   U5469 : NAND2_X1 port map( A1 => n12127, A2 => n14482, ZN => n12128);
   U5470 : NAND2_X1 port map( A1 => n12129, A2 => n12128, ZN => n12130);
   U5471 : NAND2_X1 port map( A1 => n13920, A2 => n13262, ZN => n12133);
   U5472 : NAND2_X1 port map( A1 => n14728, A2 => n14467, ZN => n12132);
   U5473 : MUX2_X1 port map( A => n14833, B => n12783, S => n12246, Z => n12137
                           );
   U5474 : NAND2_X1 port map( A1 => n14727, A2 => n12135, ZN => n12136);
   U5475 : OAI21_X1 port map( B1 => n10644, B2 => n13035, A => n12138, ZN => 
                           n12140);
   U5476 : NAND2_X1 port map( A1 => n10644, A2 => n10698, ZN => n12139);
   U5477 : NAND2_X1 port map( A1 => n12140, A2 => n12139, ZN => n13049);
   U5478 : INV_X1 port map( A => n13049, ZN => n12155);
   U5479 : MUX2_X1 port map( A => n14779, B => n14456, S => n10841, Z => n12141
                           );
   U5480 : NAND2_X1 port map( A1 => n12141, A2 => n14017, ZN => n13038);
   U5481 : MUX2_X1 port map( A => n12142, B => n10745, S => n12743, Z => n12145
                           );
   U5482 : XNOR2_X1 port map( A => n10914, B => n12671, ZN => n12143);
   U5483 : NAND2_X1 port map( A1 => n12143, A2 => n12640, ZN => n12144);
   U5484 : NAND2_X1 port map( A1 => n12145, A2 => n12144, ZN => n13037);
   U5485 : AND2_X1 port map( A1 => n13038, A2 => n13037, ZN => n12150);
   U5486 : MUX2_X1 port map( A => n14114, B => n13362, S => n8351, Z => n12148)
                           ;
   U5487 : MUX2_X1 port map( A => n12146, B => n11225, S => n12764, Z => n12147
                           );
   U5488 : OAI22_X1 port map( A1 => n12150, A2 => n12149, B1 => n13038, B2 => 
                           n13037, ZN => n13048);
   U5489 : INV_X1 port map( A => n13048, ZN => n12154);
   U5490 : NAND2_X1 port map( A1 => n12152, A2 => n12151, ZN => n13051);
   U5491 : XOR2_X1 port map( A => n12189, B => n12188, Z => n12187);
   U5492 : XNOR2_X1 port map( A => n8349, B => n8355, ZN => n12162);
   U5493 : NAND2_X1 port map( A1 => n14825, A2 => n8325, ZN => n12158);
   U5494 : OAI21_X1 port map( B1 => n8325, B2 => n14781, A => n8355, ZN => 
                           n12159);
   U5495 : NAND2_X1 port map( A1 => n12160, A2 => n12159, ZN => n12161);
   U5496 : OAI21_X1 port map( B1 => n12162, B2 => n14782, A => n12161, ZN => 
                           n13042);
   U5497 : NAND2_X1 port map( A1 => n12163, A2 => n14448, ZN => n12165);
   U5498 : NAND2_X1 port map( A1 => n14878, A2 => n8401, ZN => n12164);
   U5499 : NAND2_X1 port map( A1 => n12165, A2 => n12164, ZN => n12168);
   U5500 : XNOR2_X1 port map( A => n8352, B => n10879, ZN => n12166);
   U5501 : NAND2_X1 port map( A1 => n14789, A2 => n12166, ZN => n12167);
   U5502 : NAND2_X1 port map( A1 => n12168, A2 => n12167, ZN => n13041);
   U5503 : MUX2_X1 port map( A => n14840, B => n10645, S => n11703, Z => n12170
                           );
   U5504 : MUX2_X1 port map( A => n13442, B => n10736, S => n14451, Z => n12169
                           );
   U5505 : OAI21_X1 port map( B1 => n14121, B2 => n12170, A => n12169, ZN => 
                           n13043);
   U5506 : OAI21_X1 port map( B1 => n12172, B2 => n13043, A => n12171, ZN => 
                           n12998);
   U5507 : INV_X1 port map( A => n12998, ZN => n12185);
   U5508 : MUX2_X1 port map( A => n13347, B => n14716, S => n10742, Z => n12181
                           );
   U5509 : XNOR2_X1 port map( A => FP_A(13), B => n359, ZN => n10868);
   U5510 : NAND2_X1 port map( A1 => n12174, A2 => n12173, ZN => n12180);
   U5511 : NAND2_X1 port map( A1 => n12181, A2 => n12180, ZN => n13012);
   U5512 : NOR2_X1 port map( A1 => n14025, A2 => n13482, ZN => n13010);
   U5513 : INV_X1 port map( A => n13010, ZN => n12175);
   U5514 : NAND2_X1 port map( A1 => n12175, A2 => n11594, ZN => n12182);
   U5515 : NAND2_X1 port map( A1 => n13012, A2 => n12182, ZN => n12178);
   U5516 : MUX2_X1 port map( A => n14487, B => n13367, S => n14731, Z => n12177
                           );
   U5517 : MUX2_X1 port map( A => n13486, B => n14480, S => n13914, Z => n12176
                           );
   U5518 : NAND2_X1 port map( A1 => n13010, A2 => n14784, ZN => n12179);
   U5519 : NAND3_X1 port map( A1 => n12178, A2 => n12996, A3 => n12179, ZN => 
                           n12184);
   U5520 : AOI21_X1 port map( B1 => n12185, B2 => n12184, A => n12183, ZN => 
                           n12191);
   U5521 : INV_X1 port map( A => n12191, ZN => n12186);
   U5522 : XNOR2_X1 port map( A => n12189, B => n12188, ZN => n12190);
   U5523 : NAND2_X1 port map( A1 => n12191, A2 => n12190, ZN => n12992);
   U5524 : INV_X1 port map( A => n12992, ZN => n12192);
   U5525 : AOI21_X1 port map( B1 => n10646, B2 => n10708, A => n12192, ZN => 
                           n14824);
   U5526 : NAND2_X1 port map( A1 => n12194, A2 => n12193, ZN => n12195);
   U5527 : AND2_X1 port map( A1 => n14346, A2 => n12195, ZN => 
                           I3_SIG_out_16_port);
   U5528 : MUX2_X1 port map( A => n14020, B => n10939, S => n13450, Z => n12197
                           );
   U5529 : NAND2_X1 port map( A1 => n12230, A2 => n10726, ZN => n12196);
   U5530 : AND2_X1 port map( A1 => n12197, A2 => n12196, ZN => intadd_46_CI);
   U5531 : MUX2_X1 port map( A => n13824, B => n12163, S => n14467, Z => n12198
                           );
   U5532 : NAND2_X1 port map( A1 => n12199, A2 => n12198, ZN => n12200);
   U5533 : INV_X1 port map( A => n12200, ZN => n14111);
   U5534 : NAND2_X1 port map( A1 => n8329, A2 => n13809, ZN => n13800);
   U5535 : INV_X1 port map( A => n13800, ZN => n14109);
   U5536 : NAND2_X1 port map( A1 => n14111, A2 => n14109, ZN => n12205);
   U5537 : NAND2_X1 port map( A1 => n12200, A2 => n13800, ZN => n12203);
   U5538 : NAND2_X1 port map( A1 => n13442, A2 => n14840, ZN => n12201);
   U5539 : NAND2_X1 port map( A1 => n12201, A2 => n14460, ZN => n12202);
   U5540 : MUX2_X1 port map( A => n12202, B => n14840, S => n10841, Z => n14110
                           );
   U5541 : NAND2_X1 port map( A1 => n12203, A2 => n14110, ZN => n12204);
   U5542 : NAND2_X1 port map( A1 => n12205, A2 => n12204, ZN => n13799);
   U5543 : MUX2_X1 port map( A => n14880, B => n10886, S => n13262, Z => n12207
                           );
   U5544 : MUX2_X1 port map( A => n13819, B => n14882, S => n13823, Z => n12206
                           );
   U5545 : AND2_X1 port map( A1 => n12207, A2 => n12206, ZN => n13797);
   U5546 : OAI21_X1 port map( B1 => n13799, B2 => n14481, A => n13797, ZN => 
                           n12209);
   U5547 : NAND2_X1 port map( A1 => n13799, A2 => n14481, ZN => n12208);
   U5548 : NAND2_X1 port map( A1 => n12209, A2 => n12208, ZN => n14296);
   U5549 : XNOR2_X1 port map( A => n12211, B => n12210, ZN => n12213);
   U5550 : XNOR2_X1 port map( A => n12213, B => n12212, ZN => n12221);
   U5551 : INV_X1 port map( A => n12221, ZN => n12219);
   U5552 : MUX2_X1 port map( A => n12163, B => n14878, S => n13261, Z => n12214
                           );
   U5553 : NAND2_X1 port map( A1 => n12215, A2 => n12214, ZN => n13803);
   U5554 : NAND2_X1 port map( A1 => n10631, A2 => n14718, ZN => n13801);
   U5555 : NAND2_X1 port map( A1 => n13800, A2 => n13801, ZN => n12217);
   U5556 : NOR2_X1 port map( A1 => n13800, A2 => n13801, ZN => n12216);
   U5557 : AOI21_X1 port map( B1 => n13803, B2 => n12217, A => n12216, ZN => 
                           n12220);
   U5558 : INV_X1 port map( A => n12220, ZN => n12218);
   U5559 : NAND2_X1 port map( A1 => n12219, A2 => n12218, ZN => n14293);
   U5560 : NAND2_X1 port map( A1 => n14296, A2 => n14293, ZN => n12222);
   U5561 : NAND2_X1 port map( A1 => n12221, A2 => n12220, ZN => n14294);
   U5562 : NAND2_X1 port map( A1 => n12222, A2 => n14294, ZN => n14358);
   U5563 : XNOR2_X1 port map( A => n12224, B => n12223, ZN => n12225);
   U5564 : XNOR2_X1 port map( A => n12226, B => n12225, ZN => n14356);
   U5565 : NAND2_X1 port map( A1 => n14358, A2 => n14356, ZN => n14913);
   U5566 : MUX2_X1 port map( A => n11957, B => n11043, S => n14593, Z => n12229
                           );
   U5567 : MUX2_X1 port map( A => n10725, B => n11834, S => n14447, Z => n12228
                           );
   U5568 : NAND2_X1 port map( A1 => n12229, A2 => n12228, ZN => n12835);
   U5569 : MUX2_X1 port map( A => n14020, B => n10939, S => n12764, Z => n12232
                           );
   U5570 : NAND2_X1 port map( A1 => n12230, A2 => n14819, ZN => n12231);
   U5571 : NAND2_X1 port map( A1 => n12232, A2 => n12231, ZN => n12834);
   U5572 : AND2_X1 port map( A1 => n12835, A2 => n12834, ZN => 
                           intadd_58_A_1_port);
   U5573 : XNOR2_X1 port map( A => n12233, B => n14062, ZN => n14774);
   U5574 : INV_X1 port map( A => n14309, ZN => n12236);
   U5575 : XNOR2_X1 port map( A => n14883, B => n10841, ZN => n12234);
   U5576 : NAND2_X1 port map( A1 => n12234, A2 => n10702, ZN => n14308);
   U5577 : INV_X1 port map( A => n14308, ZN => n12235);
   U5578 : NAND2_X1 port map( A1 => n12236, A2 => n12235, ZN => n14887);
   U5579 : INV_X1 port map( A => n14887, ZN => n14888);
   U5580 : NAND2_X1 port map( A1 => EXP_out_round_2_port, A2 => 
                           EXP_out_round_3_port, ZN => n12237);
   U5581 : INV_X1 port map( A => n14435, ZN => n14929);
   U5582 : NOR2_X1 port map( A1 => n10831, A2 => n13482, ZN => 
                           intadd_62_A_0_port);
   U5583 : MUX2_X1 port map( A => n14878, B => n12163, S => n10726, Z => n12238
                           );
   U5584 : AND2_X1 port map( A1 => n12239, A2 => n12238, ZN => n14266);
   U5585 : MUX2_X1 port map( A => n13817, B => n10885, S => n11649, Z => n12241
                           );
   U5586 : MUX2_X1 port map( A => n13819, B => n14882, S => n13813, Z => n12240
                           );
   U5587 : AND2_X1 port map( A1 => n12241, A2 => n12240, ZN => n14265);
   U5588 : MUX2_X1 port map( A => n14840, B => n10645, S => n8334, Z => n12245)
                           ;
   U5589 : MUX2_X1 port map( A => n13442, B => n10738, S => n14458, Z => n12244
                           );
   U5590 : OAI21_X1 port map( B1 => n14121, B2 => n12245, A => n12244, ZN => 
                           n14123);
   U5591 : NAND2_X1 port map( A1 => n12246, A2 => n10702, ZN => n12247);
   U5592 : NAND2_X1 port map( A1 => n14449, A2 => n10702, ZN => n12674);
   U5593 : NOR2_X1 port map( A1 => n12247, A2 => n12674, ZN => n14124);
   U5594 : NAND2_X1 port map( A1 => n12247, A2 => n12674, ZN => n14125);
   U5595 : OAI21_X1 port map( B1 => n14123, B2 => n14124, A => n14125, ZN => 
                           n14264);
   U5596 : INV_X1 port map( A => intadd_61_n7, ZN => intadd_61_n1);
   U5597 : OR2_X1 port map( A1 => n12250, A2 => n12249, ZN => n12251);
   U5598 : AND2_X1 port map( A1 => n12248, A2 => n12251, ZN => 
                           I3_SIG_out_10_port);
   U5599 : NAND2_X1 port map( A1 => n12253, A2 => n14895, ZN => n12254);
   U5600 : AND2_X1 port map( A1 => n12252, A2 => n12254, ZN => 
                           I3_SIG_out_5_port);
   U5601 : AND2_X1 port map( A1 => B_EXP_7_port, A2 => A_EXP_7_port, ZN => 
                           I2_EXP_pos_int);
   U5602 : AND2_X1 port map( A1 => A_EXP_0_port, A2 => B_EXP_0_port, ZN => 
                           n12255);
   U5603 : NOR2_X1 port map( A1 => A_EXP_0_port, A2 => B_EXP_0_port, ZN => 
                           n14407);
   U5604 : OR2_X1 port map( A1 => n12255, A2 => n14407, ZN => 
                           I2_mw_I4sum_0_port);
   U5605 : NAND2_X1 port map( A1 => n14502, A2 => SIG_in_27_port, ZN => n14413)
                           ;
   U5606 : NOR2_X1 port map( A1 => n14413, A2 => n2577, ZN => n14415);
   U5607 : NAND2_X1 port map( A1 => n14415, A2 => EXP_in_2_port, ZN => n14412);
   U5608 : OR2_X1 port map( A1 => n14415, A2 => EXP_in_2_port, ZN => n12256);
   U5609 : AND2_X1 port map( A1 => n14412, A2 => n12256, ZN => 
                           I3_EXP_out_2_port);
   U5610 : NOR2_X1 port map( A1 => n14412, A2 => n14511, ZN => n12257);
   U5611 : NAND2_X1 port map( A1 => n12257, A2 => n14494, ZN => n14416);
   U5612 : OR2_X1 port map( A1 => n12257, A2 => n14494, ZN => n12258);
   U5613 : AND2_X1 port map( A1 => n14416, A2 => n12258, ZN => 
                           I3_EXP_out_4_port);
   U5614 : NAND2_X1 port map( A1 => n12260, A2 => n12259, ZN => n12262);
   U5615 : NAND2_X1 port map( A1 => n12262, A2 => n12261, ZN => n12990);
   U5616 : INV_X1 port map( A => n12990, ZN => n14765);
   U5617 : XOR2_X1 port map( A => n12265, B => n14682, Z => n14461);
   U5618 : OR2_X1 port map( A1 => n10809, A2 => n10787, ZN => n12264);
   U5619 : NAND2_X1 port map( A1 => n12265, A2 => n12264, ZN => n14485);
   U5620 : NAND2_X1 port map( A1 => n10811, A2 => n14678, ZN => n14486);
   U5621 : MUX2_X1 port map( A => n11957, B => n11043, S => n14945, Z => n12268
                           );
   U5622 : MUX2_X1 port map( A => n10725, B => n11834, S => n10743, Z => n12267
                           );
   U5623 : AND2_X1 port map( A1 => n12268, A2 => n12267, ZN => n14489);
   U5624 : XNOR2_X1 port map( A => n10823, B => n10749, ZN => n12269);
   U5625 : NAND2_X1 port map( A1 => n14776, A2 => n10765, ZN => n12271);
   U5626 : OR2_X1 port map( A1 => n10820, A2 => n10813, ZN => n12270);
   U5627 : NAND2_X1 port map( A1 => n12271, A2 => n12270, ZN => n12460);
   U5628 : NAND2_X1 port map( A1 => n12322, A2 => n12460, ZN => n12453);
   U5629 : XNOR2_X1 port map( A => n14772, B => n10813, ZN => n12448);
   U5630 : FA_X1 port map( A => n14630, B => n14629, CI => n14628, CO => n12449
                           , S => n_1339);
   U5631 : NAND2_X1 port map( A1 => n12448, A2 => n12449, ZN => n12319);
   U5632 : AND2_X1 port map( A1 => n12453, A2 => n12319, ZN => n12357);
   U5633 : INV_X1 port map( A => intadd_46_n1, ZN => n12272);
   U5634 : XNOR2_X1 port map( A => n14805, B => n14804, ZN => n12483);
   U5635 : NAND2_X1 port map( A1 => n12272, A2 => n12483, ZN => n12514);
   U5636 : NAND3_X1 port map( A1 => n10815, A2 => n10816, A3 => n14549, ZN => 
                           n12273);
   U5637 : NAND2_X1 port map( A1 => n10814, A2 => n12273, ZN => n12274);
   U5638 : NAND2_X1 port map( A1 => n10775, A2 => n12274, ZN => n12275);
   U5639 : XNOR2_X1 port map( A => n14562, B => n14561, ZN => n12296);
   U5640 : NAND2_X1 port map( A1 => n12296, A2 => n10752, ZN => n12298);
   U5641 : AND2_X1 port map( A1 => n14527, A2 => n14526, ZN => n12292);
   U5642 : NAND2_X1 port map( A1 => n14768, A2 => n12292, ZN => n12290);
   U5643 : AND3_X1 port map( A1 => n12275, A2 => n12298, A3 => n12290, ZN => 
                           n12288);
   U5644 : AOI211_X1 port map( C1 => n10776, C2 => n10814, A => n14744, B => 
                           n14743, ZN => n12281);
   U5645 : OAI21_X1 port map( B1 => n14617, B2 => n14616, A => n14615, ZN => 
                           n12278);
   U5646 : NOR2_X1 port map( A1 => n14749, A2 => n14528, ZN => n12277);
   U5647 : AOI21_X1 port map( B1 => n14564, B2 => n14563, A => n14750, ZN => 
                           n12276);
   U5648 : AOI21_X1 port map( B1 => n12278, B2 => n12277, A => n12276, ZN => 
                           n12280);
   U5649 : NAND2_X1 port map( A1 => n10632, A2 => n10643, ZN => n12279);
   U5650 : NAND4_X1 port map( A1 => n12281, A2 => n12280, A3 => n14753, A4 => 
                           n12279, ZN => n12287);
   U5651 : NAND3_X1 port map( A1 => n14753, A2 => n10816, A3 => n10815, ZN => 
                           n12282);
   U5652 : OAI21_X1 port map( B1 => n10750, B2 => n10748, A => n12282, ZN => 
                           n12284);
   U5653 : NAND2_X1 port map( A1 => n10814, A2 => n14568, ZN => n12283);
   U5654 : NAND2_X1 port map( A1 => n12284, A2 => n12283, ZN => n12286);
   U5655 : XNOR2_X1 port map( A => n14578, B => n14577, ZN => n12289);
   U5656 : NAND2_X1 port map( A1 => n14610, A2 => n12289, ZN => n12285);
   U5657 : NAND4_X1 port map( A1 => n12288, A2 => n12287, A3 => n12286, A4 => 
                           n12285, ZN => n12318);
   U5658 : INV_X1 port map( A => n12289, ZN => n12291);
   U5660 : INV_X1 port map( A => n12292, ZN => n12293);
   U5661 : NAND2_X1 port map( A1 => n14518, A2 => n12293, ZN => n12294);
   U5662 : NAND2_X1 port map( A1 => n12295, A2 => n12294, ZN => n12299);
   U5663 : INV_X1 port map( A => n12296, ZN => n12297);
   U5664 : AOI22_X1 port map( A1 => n12299, A2 => n12298, B1 => n12297, B2 => 
                           n10751, ZN => n12317);
   U5665 : INV_X1 port map( A => n12448, ZN => n12301);
   U5666 : INV_X1 port map( A => n12449, ZN => n12300);
   U5667 : NAND2_X1 port map( A1 => n12301, A2 => n12300, ZN => n12320);
   U5668 : NAND3_X1 port map( A1 => n12318, A2 => n12317, A3 => n12320, ZN => 
                           n12356);
   U5669 : AOI21_X1 port map( B1 => n10823, B2 => n10778, A => n14634, ZN => 
                           n12304);
   U5670 : INV_X1 port map( A => n12304, ZN => n12461);
   U5671 : OR2_X1 port map( A1 => n12461, A2 => intadd_46_SUM_4_port, ZN => 
                           n12355);
   U5672 : NAND4_X1 port map( A1 => n12356, A2 => n12514, A3 => n12357, A4 => 
                           n12355, ZN => n13772);
   U5673 : NOR2_X1 port map( A1 => n14625, A2 => n10777, ZN => n12302);
   U5674 : NAND2_X1 port map( A1 => n14570, A2 => n14569, ZN => n12303);
   U5675 : NAND4_X1 port map( A1 => n12302, A2 => n10823, A3 => n10749, A4 => 
                           n12303, ZN => n12359);
   U5676 : INV_X1 port map( A => n12359, ZN => n12306);
   U5677 : OAI211_X1 port map( C1 => n10823, C2 => n10778, A => n12303, B => 
                           n14644, ZN => n12305);
   U5678 : NAND2_X1 port map( A1 => n12305, A2 => n12304, ZN => n12358);
   U5679 : OAI211_X1 port map( C1 => n10853, C2 => n12306, A => n12514, B => 
                           n12358, ZN => n13768);
   U5680 : INV_X1 port map( A => n12483, ZN => n12307);
   U5681 : NAND2_X1 port map( A1 => intadd_46_n1, A2 => n12307, ZN => n13765);
   U5682 : NAND2_X1 port map( A1 => n13768, A2 => n13765, ZN => n12570);
   U5683 : INV_X1 port map( A => n12570, ZN => n12308);
   U5684 : NAND2_X1 port map( A1 => n13772, A2 => n12308, ZN => n14321);
   U5685 : XNOR2_X1 port map( A => n14633, B => n14632, ZN => n12310);
   U5686 : XNOR2_X1 port map( A => n10780, B => n14573, ZN => n12309);
   U5687 : XNOR2_X1 port map( A => n12310, B => n12309, ZN => n12373);
   U5688 : OAI21_X1 port map( B1 => n14804, B2 => n10768, A => n10764, ZN => 
                           n12312);
   U5689 : NAND2_X1 port map( A1 => n14804, A2 => n10768, ZN => n12311);
   U5690 : NAND2_X1 port map( A1 => n12312, A2 => n12311, ZN => n12372);
   U5691 : OR2_X1 port map( A1 => n12373, A2 => n12372, ZN => n14319);
   U5692 : NAND2_X1 port map( A1 => n12373, A2 => n12372, ZN => n14318);
   U5693 : AOI21_X1 port map( B1 => n14321, B2 => n14319, A => n12517, ZN => 
                           n12316);
   U5694 : XNOR2_X1 port map( A => n14550, B => n10779, ZN => n12313);
   U5695 : XNOR2_X1 port map( A => n12313, B => n14655, ZN => n12374);
   U5696 : NAND2_X1 port map( A1 => n14599, A2 => n14598, ZN => n12314);
   U5697 : NAND2_X1 port map( A1 => n12314, A2 => n14831, ZN => n12371);
   U5698 : OR2_X1 port map( A1 => n12374, A2 => n12371, ZN => n12516);
   U5699 : NAND2_X1 port map( A1 => n12374, A2 => n12371, ZN => n12324);
   U5700 : NAND2_X1 port map( A1 => n12516, A2 => n12324, ZN => n12315);
   U5701 : XNOR2_X1 port map( A => n12316, B => n12315, ZN => n14490);
   U5702 : NAND2_X1 port map( A1 => n12318, A2 => n12317, ZN => n12451);
   U5703 : NAND2_X1 port map( A1 => n12451, A2 => n12319, ZN => n12321);
   U5704 : NAND2_X1 port map( A1 => n12321, A2 => n12320, ZN => n12470);
   U5705 : INV_X1 port map( A => n12460, ZN => n12455);
   U5706 : XNOR2_X1 port map( A => n12322, B => n12455, ZN => n12323);
   U5707 : XOR2_X1 port map( A => n12470, B => n12323, Z => n14491);
   U5708 : INV_X1 port map( A => n12513, ZN => n12548);
   U5709 : AOI21_X1 port map( B1 => n12516, B2 => n12517, A => n12518, ZN => 
                           n12551);
   U5710 : INV_X1 port map( A => n12551, ZN => n12325);
   U5711 : AOI21_X1 port map( B1 => n14321, B2 => n12513, A => n12325, ZN => 
                           n12332);
   U5712 : NAND2_X1 port map( A1 => n14535, A2 => n14534, ZN => n12364);
   U5713 : NAND2_X1 port map( A1 => n14823, A2 => n12364, ZN => n12326);
   U5714 : XNOR2_X1 port map( A => n12326, B => n14657, ZN => n12330);
   U5715 : XNOR2_X1 port map( A => n10779, B => n14560, ZN => n12327);
   U5716 : NAND2_X1 port map( A1 => n12327, A2 => n14638, ZN => n12328);
   U5717 : NAND2_X1 port map( A1 => n12328, A2 => n14654, ZN => n12329);
   U5718 : NOR2_X1 port map( A1 => n12330, A2 => n12329, ZN => n12550);
   U5719 : INV_X1 port map( A => n12550, ZN => n12376);
   U5720 : NAND2_X1 port map( A1 => n12330, A2 => n12329, ZN => n12549);
   U5721 : NAND2_X1 port map( A1 => n12376, A2 => n12549, ZN => n12331);
   U5722 : XNOR2_X1 port map( A => n12332, B => n12331, ZN => n14517);
   U5723 : XNOR2_X1 port map( A => n12252, B => n14495, ZN => I3_SIG_out_6_port
                           );
   U5724 : INV_X1 port map( A => FP_A(12), ZN => n12333);
   U5725 : NOR2_X1 port map( A1 => FP_A(13), A2 => n12333, ZN => n14582);
   U5726 : NAND2_X1 port map( A1 => n14582, A2 => FP_A(11), ZN => n14583);
   U5727 : NAND2_X1 port map( A1 => n14922, A2 => n10807, ZN => FP_Z(22));
   U5728 : NAND2_X1 port map( A1 => n12068, A2 => FP_A(7), ZN => n14595);
   U5729 : NAND2_X1 port map( A1 => n12334, A2 => FP_A(3), ZN => n14603);
   U5730 : NAND2_X1 port map( A1 => n14603, A2 => n14591, ZN => n14592);
   U5731 : NAND2_X1 port map( A1 => n14609, A2 => n10807, ZN => n12692);
   U5732 : INV_X1 port map( A => n12692, ZN => n12478);
   U5733 : OAI211_X1 port map( C1 => n14576, C2 => n14575, A => n10812, B => 
                           n14574, ZN => n12335);
   U5734 : NAND2_X1 port map( A1 => n12478, A2 => n12335, ZN => FP_Z(27));
   U5735 : NAND2_X1 port map( A1 => n12478, A2 => n14930, ZN => FP_Z(29));
   U5736 : NAND2_X1 port map( A1 => n12478, A2 => n10826, ZN => FP_Z(28));
   U5737 : NOR2_X1 port map( A1 => n8379, A2 => n2579, ZN => n12352);
   U5738 : NAND2_X1 port map( A1 => n14436, A2 => n12352, ZN => n14441);
   U5739 : NAND4_X1 port map( A1 => n10970, A2 => n14485, A3 => n14461, A4 => 
                           n2563, ZN => n12337);
   U5740 : NAND4_X1 port map( A1 => n14462, A2 => n14486, A3 => n2573, A4 => 
                           n2562, ZN => n12336);
   U5741 : NOR2_X1 port map( A1 => n12337, A2 => n12336, ZN => n12341);
   U5742 : NAND4_X1 port map( A1 => n2574, A2 => n2560, A3 => n2572, A4 => 
                           n2561, ZN => n12339);
   U5743 : NAND4_X1 port map( A1 => n2570, A2 => n2559, A3 => n2571, A4 => 
                           n2557, ZN => n12338);
   U5744 : NOR2_X1 port map( A1 => n12339, A2 => n12338, ZN => n12340);
   U5745 : NAND2_X1 port map( A1 => n12341, A2 => n12340, ZN => n12348);
   U5746 : AND4_X1 port map( A1 => n2569, A2 => n2558, A3 => n2556, A4 => n2568
                           , ZN => n12346);
   U5747 : OAI211_X1 port map( C1 => n12342, C2 => n14687, A => n14686, B => 
                           n14685, ZN => n12343);
   U5748 : NAND2_X1 port map( A1 => n2587, A2 => n14446, ZN => n12344);
   U5749 : NOR2_X1 port map( A1 => n12343, A2 => n12344, ZN => n12345);
   U5750 : NAND4_X1 port map( A1 => n12346, A2 => n12345, A3 => n2565, A4 => 
                           n14921, ZN => n12347);
   U5751 : OAI21_X1 port map( B1 => n12348, B2 => n12347, A => n2611, ZN => 
                           n12349);
   U5752 : AND2_X1 port map( A1 => n14446, A2 => n2584, ZN => n12350);
   U5753 : NOR2_X1 port map( A1 => n14924, A2 => n12350, ZN => n14432);
   U5754 : AND4_X1 port map( A1 => EXP_out_round_7_port, A2 => 
                           EXP_out_round_4_port, A3 => EXP_out_round_1_port, A4
                           => EXP_out_round_3_port, ZN => n12351);
   U5755 : NAND4_X1 port map( A1 => n14432, A2 => EXP_out_round_2_port, A3 => 
                           n12352, A4 => n12351, ZN => n12353);
   U5756 : AND2_X1 port map( A1 => n12353, A2 => n8385, ZN => n12354);
   U5757 : OAI21_X1 port map( B1 => n10681, B2 => n2613, A => n12354, ZN => 
                           n14428);
   U5758 : NAND2_X1 port map( A1 => n10937, A2 => n14428, ZN => n14919);
   U5759 : OR2_X1 port map( A1 => n12692, A2 => n14642, ZN => FP_Z(23));
   U5760 : OR2_X1 port map( A1 => n12692, A2 => n14643, ZN => FP_Z(25));
   U5761 : OR2_X1 port map( A1 => n12692, A2 => n14927, ZN => FP_Z(26));
   U5762 : NAND3_X1 port map( A1 => n12357, A2 => n12356, A3 => n12355, ZN => 
                           n12482);
   U5763 : NAND2_X1 port map( A1 => intadd_46_SUM_4_port, A2 => n12358, ZN => 
                           n12360);
   U5764 : NAND2_X1 port map( A1 => n12360, A2 => n12359, ZN => n12480);
   U5765 : INV_X1 port map( A => n13765, ZN => n12361);
   U5766 : NOR2_X1 port map( A1 => n12480, A2 => n12361, ZN => n12362);
   U5767 : NAND2_X1 port map( A1 => n12482, A2 => n12362, ZN => n12564);
   U5768 : XNOR2_X1 port map( A => n14548, B => n14547, ZN => n12368);
   U5769 : XNOR2_X1 port map( A => n14530, B => n14529, ZN => n12363);
   U5770 : XNOR2_X1 port map( A => n12368, B => n12363, ZN => n12377);
   U5771 : NAND2_X1 port map( A1 => n14823, A2 => n14559, ZN => n12366);
   U5772 : NAND2_X1 port map( A1 => n14823, A2 => n14558, ZN => n12365);
   U5773 : NAND3_X1 port map( A1 => n12366, A2 => n12365, A3 => n12364, ZN => 
                           n12378);
   U5774 : NOR2_X1 port map( A1 => n12377, A2 => n12378, ZN => n12557);
   U5775 : XNOR2_X1 port map( A => n10772, B => n14590, ZN => n12367);
   U5776 : XNOR2_X1 port map( A => n12367, B => n14645, ZN => n12524);
   U5777 : INV_X1 port map( A => n12524, ZN => n12379);
   U5778 : INV_X1 port map( A => n12368, ZN => n12369);
   U5779 : NAND2_X1 port map( A1 => n12369, A2 => n14631, ZN => n12370);
   U5780 : NAND2_X1 port map( A1 => n12370, A2 => n14651, ZN => n12523);
   U5781 : INV_X1 port map( A => n12523, ZN => n12380);
   U5782 : NAND2_X1 port map( A1 => n12379, A2 => n12380, ZN => n12575);
   U5783 : AND4_X2 port map( A1 => n12513, A2 => n12519, A3 => n12575, A4 => 
                           n12514, ZN => n12563);
   U5784 : NAND2_X1 port map( A1 => n12564, A2 => n12563, ZN => n13702);
   U5785 : AND2_X1 port map( A1 => n12374, A2 => n12371, ZN => n12518);
   U5786 : AND2_X1 port map( A1 => n12373, A2 => n12372, ZN => n12517);
   U5787 : OR2_X1 port map( A1 => n12374, A2 => n14522, ZN => n12375);
   U5788 : OAI211_X1 port map( C1 => n12518, C2 => n12517, A => n12376, B => 
                           n12375, ZN => n12384);
   U5789 : NAND2_X1 port map( A1 => n12377, A2 => n12378, ZN => n12555);
   U5790 : AND2_X1 port map( A1 => n12549, A2 => n12555, ZN => n13767);
   U5791 : NAND2_X1 port map( A1 => n12524, A2 => n12523, ZN => n12568);
   U5792 : AND2_X1 port map( A1 => n13767, A2 => n12568, ZN => n12383);
   U5793 : INV_X1 port map( A => n12557, ZN => n12520);
   U5794 : OAI21_X1 port map( B1 => n12557, B2 => n12380, A => n12379, ZN => 
                           n12381);
   U5795 : OAI21_X1 port map( B1 => n12520, B2 => n12523, A => n12381, ZN => 
                           n12382);
   U5796 : AOI21_X1 port map( B1 => n12384, B2 => n12383, A => n12382, ZN => 
                           n12502);
   U5797 : XNOR2_X1 port map( A => n14627, B => n10770, ZN => n14333);
   U5798 : FA_X1 port map( A => n10781, B => n14637, CI => n14636, CO => n14334
                           , S => n_1340);
   U5799 : AND2_X1 port map( A1 => n14333, A2 => n14334, ZN => n12580);
   U5801 : INV_X1 port map( A => n12388, ZN => n12386);
   U5802 : XNOR2_X1 port map( A => n14842, B => n14587, ZN => n12387);
   U5803 : INV_X1 port map( A => n12387, ZN => n12385);
   U5806 : NAND2_X1 port map( A1 => n12388, A2 => n12387, ZN => n13608);
   U5807 : XNOR2_X1 port map( A => n14588, B => n10782, ZN => n13604);
   U5808 : INV_X1 port map( A => n13604, ZN => n12390);
   U5809 : AND2_X1 port map( A1 => n14554, A2 => n10769, ZN => n13605);
   U5810 : INV_X1 port map( A => n13605, ZN => n12389);
   U5811 : NAND2_X1 port map( A1 => n12390, A2 => n12389, ZN => n12391);
   U5812 : NAND2_X1 port map( A1 => n13608, A2 => n12391, ZN => n12407);
   U5813 : NOR2_X1 port map( A1 => n13607, A2 => n12407, ZN => n12611);
   U5814 : FA_X1 port map( A => n10773, B => n14659, CI => n10771, CO => n12419
                           , S => n_1341);
   U5815 : XNOR2_X1 port map( A => n10781, B => n14537, ZN => n12392);
   U5816 : XOR2_X1 port map( A => n12392, B => n14650, Z => n12420);
   U5817 : OR2_X1 port map( A1 => n12419, A2 => n12420, ZN => n12606);
   U5818 : XNOR2_X1 port map( A => n14539, B => n14538, ZN => n13785);
   U5819 : NAND2_X1 port map( A1 => n14589, A2 => n10783, ZN => n13786);
   U5820 : NOR2_X1 port map( A1 => n13785, A2 => n13786, ZN => n13757);
   U5821 : NOR2_X1 port map( A1 => n13757, A2 => n12425, ZN => n12421);
   U5822 : FA_X1 port map( A => n14612, B => n14611, CI => n10782, CO => n12406
                           , S => n_1342);
   U5823 : INV_X1 port map( A => n12406, ZN => n12394);
   U5824 : XNOR2_X1 port map( A => n14614, B => n14613, ZN => n12405);
   U5825 : INV_X1 port map( A => n12405, ZN => n12393);
   U5826 : NAND2_X1 port map( A1 => n12394, A2 => n12393, ZN => n12617);
   U5827 : AND3_X1 port map( A1 => n12606, A2 => n12421, A3 => n12617, ZN => 
                           n12409);
   U5828 : XNOR2_X1 port map( A => n10784, B => n10785, ZN => n12395);
   U5829 : XNOR2_X1 port map( A => n14556, B => n14555, ZN => n12397);
   U5830 : INV_X1 port map( A => n12397, ZN => n12398);
   U5831 : XNOR2_X1 port map( A => n12395, B => n12398, ZN => n12494);
   U5832 : INV_X1 port map( A => n12494, ZN => n12411);
   U5833 : NAND2_X1 port map( A1 => n10754, A2 => n14626, ZN => n12396);
   U5834 : AOI22_X1 port map( A1 => n12396, A2 => n10772, B1 => n10753, B2 => 
                           n14656, ZN => n12493);
   U5835 : INV_X1 port map( A => n12493, ZN => n12404);
   U5836 : NAND2_X1 port map( A1 => n12411, A2 => n12404, ZN => n12603);
   U5837 : NAND2_X1 port map( A1 => n12397, A2 => n10785, ZN => n12399);
   U5838 : INV_X1 port map( A => n12607, ZN => n12402);
   U5839 : XNOR2_X1 port map( A => n10771, B => n14552, ZN => n12400);
   U5840 : XNOR2_X1 port map( A => n12400, B => n10774, ZN => n12605);
   U5841 : INV_X1 port map( A => n12605, ZN => n12403);
   U5842 : NAND4_X1 port map( A1 => n12409, A2 => n12611, A3 => n12603, A4 => 
                           n12578, ZN => n12401);
   U5843 : NOR2_X1 port map( A1 => n12502, A2 => n12401, ZN => n13701);
   U5844 : NAND2_X1 port map( A1 => n13701, A2 => n13702, ZN => n13731);
   U5845 : OAI21_X1 port map( B1 => n12404, B2 => n12403, A => n12402, ZN => 
                           n12408);
   U5846 : NAND2_X1 port map( A1 => n13605, A2 => n13604, ZN => n12612);
   U5847 : NAND2_X1 port map( A1 => n12406, A2 => n12405, ZN => n12616);
   U5848 : AND2_X1 port map( A1 => n12612, A2 => n12616, ZN => n13762);
   U5849 : NAND2_X1 port map( A1 => n12407, A2 => n13762, ZN => n12416);
   U5850 : AND2_X1 port map( A1 => n12408, A2 => n12416, ZN => n12415);
   U5851 : INV_X1 port map( A => n13607, ZN => n12410);
   U5852 : OR2_X1 port map( A1 => n12493, A2 => n12605, ZN => n12413);
   U5853 : NAND2_X1 port map( A1 => n12607, A2 => n12605, ZN => n12577);
   U5854 : NAND2_X1 port map( A1 => n12411, A2 => n12577, ZN => n12412);
   U5856 : AND2_X1 port map( A1 => n12416, A2 => n12617, ZN => n12587);
   U5857 : NAND2_X1 port map( A1 => n13607, A2 => n13762, ZN => n12588);
   U5858 : INV_X1 port map( A => n14333, ZN => n12418);
   U5859 : INV_X1 port map( A => n14334, ZN => n12417);
   U5860 : NAND2_X1 port map( A1 => n12418, A2 => n12417, ZN => n12585);
   U5861 : NAND2_X1 port map( A1 => n12420, A2 => n12419, ZN => n13776);
   U5862 : NAND4_X1 port map( A1 => n12597, A2 => n13762, A3 => n12585, A4 => 
                           n13776, ZN => n13761);
   U5863 : NAND4_X1 port map( A1 => n12587, A2 => n12588, A3 => n12421, A4 => 
                           n13761, ZN => n13686);
   U5864 : NAND2_X1 port map( A1 => n10783, A2 => n14546, ZN => n12422);
   U5865 : AND2_X1 port map( A1 => n12422, A2 => n14618, ZN => n13788);
   U5866 : NAND2_X1 port map( A1 => n13788, A2 => n13785, ZN => n13758);
   U5867 : OR2_X1 port map( A1 => n10817, A2 => n12423, ZN => n12424);
   U5868 : NAND2_X1 port map( A1 => n13758, A2 => n12424, ZN => n12427);
   U5869 : INV_X1 port map( A => n12425, ZN => n12426);
   U5870 : NAND2_X1 port map( A1 => n12427, A2 => n12426, ZN => n13682);
   U5871 : NAND2_X1 port map( A1 => n10824, A2 => n10822, ZN => n13709);
   U5872 : OAI21_X1 port map( B1 => n14533, B2 => n14532, A => n14531, ZN => 
                           n12531);
   U5873 : NAND2_X1 port map( A1 => n10819, A2 => n12531, ZN => n12538);
   U5874 : NAND2_X1 port map( A1 => n13709, A2 => n12538, ZN => n14365);
   U5875 : XNOR2_X1 port map( A => n14623, B => n14622, ZN => n13729);
   U5876 : NAND2_X1 port map( A1 => n10786, A2 => n14551, ZN => n12428);
   U5877 : NAND2_X1 port map( A1 => n12428, A2 => n14624, ZN => n12431);
   U5878 : AND2_X1 port map( A1 => n13729, A2 => n12431, ZN => n12429);
   U5879 : NOR2_X1 port map( A1 => n14365, A2 => n12429, ZN => n12430);
   U5880 : XNOR2_X1 port map( A => n14608, B => n10786, ZN => n13743);
   U5881 : FA_X1 port map( A => n14544, B => n14543, CI => n14542, CO => n12529
                           , S => n12423);
   U5882 : NAND2_X1 port map( A1 => n13743, A2 => n12529, ZN => n13732);
   U5883 : NAND2_X1 port map( A1 => n12430, A2 => n13732, ZN => n14364);
   U5884 : NAND2_X1 port map( A1 => n12528, A2 => n13749, ZN => n12440);
   U5885 : INV_X1 port map( A => n13729, ZN => n12432);
   U5886 : INV_X1 port map( A => n13743, ZN => n12433);
   U5887 : INV_X1 port map( A => n12529, ZN => n13742);
   U5888 : NAND3_X1 port map( A1 => n12432, A2 => n12433, A3 => n13742, ZN => 
                           n12435);
   U5889 : INV_X1 port map( A => n12431, ZN => n13730);
   U5890 : NAND2_X1 port map( A1 => n12432, A2 => n13730, ZN => n12530);
   U5891 : NAND3_X1 port map( A1 => n12433, A2 => n13730, A3 => n13742, ZN => 
                           n12434);
   U5892 : NAND4_X1 port map( A1 => n12435, A2 => n12530, A3 => n12434, A4 => 
                           n13690, ZN => n14368);
   U5893 : NOR2_X1 port map( A1 => n10824, A2 => n10822, ZN => n14366);
   U5894 : INV_X1 port map( A => n12538, ZN => n13689);
   U5895 : AOI21_X1 port map( B1 => n13689, B2 => n10822, A => n10818, ZN => 
                           n12438);
   U5896 : NAND2_X1 port map( A1 => n12538, A2 => n10821, ZN => n12436);
   U5897 : NAND2_X1 port map( A1 => n12436, A2 => n10824, ZN => n12437);
   U5898 : OAI211_X1 port map( C1 => n14368, C2 => n14366, A => n12438, B => 
                           n12437, ZN => n12439);
   U5899 : INV_X1 port map( A => n13749, ZN => n12441);
   U5900 : NOR2_X1 port map( A1 => n12441, A2 => n14689, ZN => n12445);
   U5901 : INV_X1 port map( A => n13752, ZN => n12442);
   U5902 : NAND2_X1 port map( A1 => n12442, A2 => n14694, ZN => n12443);
   U5903 : AOI21_X1 port map( B1 => n12443, B2 => n14696, A => n14695, ZN => 
                           n12444);
   U5904 : AOI21_X1 port map( B1 => n12528, B2 => n12445, A => n12444, ZN => 
                           n12446);
   U5905 : XNOR2_X1 port map( A => n2583, B => n14729, ZN => I3_EXP_out_0_port)
                           ;
   U5906 : XOR2_X1 port map( A => n12449, B => n12448, Z => n12450);
   U5907 : XOR2_X1 port map( A => n12451, B => n12450, Z => n12473);
   U5908 : XNOR2_X1 port map( A => n12304, B => n10853, ZN => n12454);
   U5909 : INV_X1 port map( A => n12454, ZN => n12452);
   U5910 : OAI21_X1 port map( B1 => n12322, B2 => n12460, A => n12452, ZN => 
                           n12471);
   U5911 : NAND3_X1 port map( A1 => n12470, A2 => n12454, A3 => n12453, ZN => 
                           n12469);
   U5912 : AND2_X1 port map( A1 => n12461, A2 => n12455, ZN => n12457);
   U5913 : OAI21_X1 port map( B1 => n12455, B2 => n12461, A => n12322, ZN => 
                           n12456);
   U5914 : OAI21_X1 port map( B1 => n12322, B2 => n12457, A => n12456, ZN => 
                           n12459);
   U5915 : INV_X1 port map( A => n10853, ZN => n12458);
   U5916 : NAND2_X1 port map( A1 => n12459, A2 => n12458, ZN => n12467);
   U5917 : NOR2_X1 port map( A1 => n12461, A2 => n12460, ZN => n12464);
   U5918 : NAND2_X1 port map( A1 => n12461, A2 => n12460, ZN => n12462);
   U5919 : NAND2_X1 port map( A1 => n12322, A2 => n12462, ZN => n12463);
   U5920 : OAI21_X1 port map( B1 => n12322, B2 => n12464, A => n12463, ZN => 
                           n12465);
   U5921 : NAND2_X1 port map( A1 => n12465, A2 => n10853, ZN => n12466);
   U5922 : NAND2_X1 port map( A1 => n12467, A2 => n12466, ZN => n12468);
   U5923 : OAI211_X1 port map( C1 => n12471, C2 => n12470, A => n12469, B => 
                           n12468, ZN => n12472);
   U5924 : INV_X1 port map( A => n12472, ZN => n12486);
   U5925 : MUX2_X1 port map( A => n12473, B => n12486, S => n14323, Z => n14697
                           );
   U5926 : NOR2_X1 port map( A1 => n14697, A2 => n14491, ZN => n14619);
   U5927 : AND2_X1 port map( A1 => n14891, A2 => n14890, ZN => n12474);
   U5928 : NOR2_X1 port map( A1 => n14894, A2 => n12474, ZN => n10596);
   U5929 : AND2_X1 port map( A1 => n10681, A2 => n14931, ZN => n14932);
   U5930 : INV_X1 port map( A => n14663, ZN => n12476);
   U5931 : NAND2_X1 port map( A1 => n12476, A2 => n13843, ZN => n14652);
   U5932 : OAI211_X1 port map( C1 => n14567, C2 => n14566, A => n10746, B => 
                           n14565, ZN => n12477);
   U5933 : NAND2_X1 port map( A1 => n12478, A2 => n12477, ZN => FP_Z(24));
   U5934 : NOR2_X1 port map( A1 => FP_A(4), A2 => n14596, ZN => n12479);
   U5935 : NAND2_X1 port map( A1 => n12479, A2 => n14541, ZN => n14540);
   U5936 : XNOR2_X1 port map( A => n14894, B => n14892, ZN => I3_SIG_out_4_port
                           );
   U5937 : INV_X1 port map( A => n12480, ZN => n12481);
   U5938 : NAND2_X1 port map( A1 => n12482, A2 => n12481, ZN => n12485);
   U5939 : XNOR2_X1 port map( A => intadd_46_n1, B => n12483, ZN => n12484);
   U5940 : XOR2_X1 port map( A => n12485, B => n12484, Z => n14322);
   U5941 : MUX2_X1 port map( A => n12486, B => n14322, S => n14323, Z => n14658
                           );
   U5942 : INV_X1 port map( A => n14658, ZN => n14545);
   U5943 : NAND3_X1 port map( A1 => FP_A(14), A2 => FP_A(13), A3 => n384, ZN =>
                           n14660);
   U5944 : NAND2_X1 port map( A1 => n14668, A2 => n14605, ZN => n14604);
   U5946 : XOR2_X1 port map( A => n14605, B => n14667, Z => n14666);
   U5947 : XNOR2_X1 port map( A => n14702, B => FP_A(3), ZN => n14606);
   U5948 : XNOR2_X1 port map( A => n14602, B => n384, ZN => n14669);
   U5949 : INV_X1 port map( A => n10936, ZN => n14920);
   U5950 : OAI22_X1 port map( A1 => n10760, A2 => n12491, B1 => n12492, B2 => 
                           n10762, ZN => FP_Z(19));
   U5951 : OAI22_X1 port map( A1 => n10805, A2 => n12490, B1 => n12489, B2 => 
                           n14680, ZN => FP_Z(0));
   U5952 : OAI22_X1 port map( A1 => n10802, A2 => n12489, B1 => n12491, B2 => 
                           n10801, ZN => FP_Z(4));
   U5953 : OAI22_X1 port map( A1 => n10805, A2 => n12489, B1 => n12490, B2 => 
                           n10804, ZN => FP_Z(1));
   U5954 : OAI22_X1 port map( A1 => n10799, A2 => n12490, B1 => n12492, B2 => 
                           n10800, ZN => FP_Z(6));
   U5955 : OAI22_X1 port map( A1 => n10795, A2 => n12491, B1 => n12489, B2 => 
                           n10796, ZN => FP_Z(10));
   U5956 : OAI22_X1 port map( A1 => n10797, A2 => n12490, B1 => n12489, B2 => 
                           n10798, ZN => FP_Z(8));
   U5957 : OAI22_X1 port map( A1 => n10763, A2 => n12491, B1 => n12492, B2 => 
                           n10790, ZN => FP_Z(16));
   U5958 : OAI22_X1 port map( A1 => n10802, A2 => n12490, B1 => n12492, B2 => 
                           n10803, ZN => FP_Z(3));
   U5959 : OAI22_X1 port map( A1 => n10794, A2 => n12489, B1 => n12491, B2 => 
                           n10793, ZN => FP_Z(12));
   U5960 : OAI22_X1 port map( A1 => n10798, A2 => n12491, B1 => n12489, B2 => 
                           n10799, ZN => FP_Z(7));
   U5961 : OAI22_X1 port map( A1 => n10794, A2 => n12490, B1 => n12489, B2 => 
                           n10795, ZN => FP_Z(11));
   U5962 : OAI22_X1 port map( A1 => n10800, A2 => n12491, B1 => n12492, B2 => 
                           n10801, ZN => FP_Z(5));
   U5963 : OAI22_X1 port map( A1 => n10797, A2 => n12492, B1 => n12490, B2 => 
                           n10796, ZN => FP_Z(9));
   U5964 : OAI22_X1 port map( A1 => n10791, A2 => n12490, B1 => n12492, B2 => 
                           n10792, ZN => FP_Z(14));
   U5965 : OAI22_X1 port map( A1 => n10803, A2 => n12491, B1 => n12489, B2 => 
                           n10804, ZN => FP_Z(2));
   U5966 : OAI22_X1 port map( A1 => n10792, A2 => n12490, B1 => n12492, B2 => 
                           n10793, ZN => FP_Z(13));
   U5967 : OAI22_X1 port map( A1 => n10761, A2 => n12491, B1 => n12489, B2 => 
                           n10763, ZN => FP_Z(17));
   U5968 : OAI22_X1 port map( A1 => n10791, A2 => n12489, B1 => n12490, B2 => 
                           n10790, ZN => FP_Z(15));
   U5969 : OAI22_X1 port map( A1 => n10761, A2 => n12492, B1 => n12491, B2 => 
                           n10762, ZN => FP_Z(18));
   U5970 : OAI22_X1 port map( A1 => n10760, A2 => n12492, B1 => n12490, B2 => 
                           n10747, ZN => FP_Z(20));
   U5971 : OAI22_X1 port map( A1 => n10747, A2 => n12492, B1 => n12491, B2 => 
                           n14681, ZN => FP_Z(21));
   U5972 : NAND2_X1 port map( A1 => n12494, A2 => n12493, ZN => n12598);
   U5973 : AND2_X1 port map( A1 => n12598, A2 => n12577, ZN => n12496);
   U5974 : AND2_X1 port map( A1 => n12606, A2 => n13776, ZN => n12495);
   U5975 : NAND2_X1 port map( A1 => n12496, A2 => n12495, ZN => n12503);
   U5976 : OR2_X1 port map( A1 => n13702, A2 => n12503, ZN => n12508);
   U5977 : INV_X1 port map( A => n12578, ZN => n12500);
   U5978 : INV_X1 port map( A => n12495, ZN => n12504);
   U5979 : INV_X1 port map( A => n12496, ZN => n12497);
   U5980 : NAND2_X1 port map( A1 => n12497, A2 => n12578, ZN => n12498);
   U5981 : NAND2_X1 port map( A1 => n12498, A2 => n12504, ZN => n12499);
   U5982 : OAI21_X1 port map( B1 => n12500, B2 => n12504, A => n12499, ZN => 
                           n12507);
   U5983 : INV_X1 port map( A => n12603, ZN => n12501);
   U5984 : NOR2_X1 port map( A1 => n10699, A2 => n12501, ZN => n12510);
   U5985 : OR2_X1 port map( A1 => n12510, A2 => n12503, ZN => n12506);
   U5986 : NAND4_X1 port map( A1 => n10728, A2 => n12510, A3 => n12578, A4 => 
                           n12504, ZN => n12505);
   U5987 : NAND4_X1 port map( A1 => n12508, A2 => n12507, A3 => n12506, A4 => 
                           n12505, ZN => I2_dtemp_33_port);
   U5988 : INV_X1 port map( A => n12598, ZN => n12509);
   U5989 : AOI21_X1 port map( B1 => n10728, B2 => n12510, A => n12509, ZN => 
                           n12512);
   U5990 : AND2_X1 port map( A1 => n12577, A2 => n12578, ZN => n12511);
   U5991 : XNOR2_X1 port map( A => n12512, B => n12511, ZN => n10593);
   U5992 : NAND2_X1 port map( A1 => n12513, A2 => n12519, ZN => n12574);
   U5993 : INV_X1 port map( A => n12514, ZN => n12515);
   U5994 : NOR2_X1 port map( A1 => n12574, A2 => n12515, ZN => n12522);
   U5995 : NAND3_X1 port map( A1 => n12519, A2 => n12517, A3 => n12516, ZN => 
                           n13769);
   U5996 : NAND2_X1 port map( A1 => n12519, A2 => n12518, ZN => n12569);
   U5997 : INV_X1 port map( A => n13767, ZN => n12521);
   U5998 : NAND2_X1 port map( A1 => n12521, A2 => n12520, ZN => n12573);
   U5999 : NAND3_X1 port map( A1 => n13769, A2 => n12569, A3 => n12573, ZN => 
                           n12560);
   U6000 : AOI21_X1 port map( B1 => n12564, B2 => n12522, A => n12560, ZN => 
                           n12527);
   U6001 : XNOR2_X1 port map( A => n12524, B => n12523, ZN => n12526);
   U6002 : NAND2_X1 port map( A1 => n12527, A2 => n12526, ZN => n12525);
   U6003 : OAI21_X1 port map( B1 => n12527, B2 => n12526, A => n12525, ZN => 
                           I2_dtemp_30_port);
   U6004 : OR2_X1 port map( A1 => n13743, A2 => n12529, ZN => n13734);
   U6005 : NAND2_X1 port map( A1 => n12530, A2 => n13734, ZN => n13685);
   U6006 : INV_X1 port map( A => n13685, ZN => n12533);
   U6007 : XNOR2_X1 port map( A => n10819, B => n12531, ZN => n12540);
   U6008 : INV_X1 port map( A => n12540, ZN => n12532);
   U6009 : NAND2_X1 port map( A1 => n12533, A2 => n12532, ZN => n12547);
   U6010 : NAND2_X1 port map( A1 => n13732, A2 => n13730, ZN => n12534);
   U6011 : NAND2_X1 port map( A1 => n12534, A2 => n13729, ZN => n12536);
   U6012 : OR2_X1 port map( A1 => n13732, A2 => n13730, ZN => n12535);
   U6013 : NAND2_X1 port map( A1 => n12536, A2 => n12535, ZN => n13691);
   U6014 : NOR2_X1 port map( A1 => n13691, A2 => n13685, ZN => n12537);
   U6015 : NAND2_X1 port map( A1 => n10700, A2 => n12537, ZN => n12543);
   U6016 : INV_X1 port map( A => n13691, ZN => n12541);
   U6017 : NAND2_X1 port map( A1 => n13690, A2 => n12538, ZN => n12539);
   U6018 : NAND2_X1 port map( A1 => n12541, A2 => n12539, ZN => n12544);
   U6019 : OAI21_X1 port map( B1 => n12541, B2 => n12540, A => n12544, ZN => 
                           n12542);
   U6020 : NAND2_X1 port map( A1 => n12543, A2 => n12542, ZN => n12546);
   U6022 : OR2_X1 port map( A1 => n13747, A2 => n12544, ZN => n12545);
   U6023 : OAI211_X1 port map( C1 => n14373, C2 => n12547, A => n12546, B => 
                           n12545, ZN => I2_dtemp_42_port);
   U6024 : NOR2_X1 port map( A1 => n12548, A2 => n12550, ZN => n12553);
   U6025 : OAI21_X1 port map( B1 => n12551, B2 => n12550, A => n12549, ZN => 
                           n12552);
   U6026 : AOI21_X1 port map( B1 => n14321, B2 => n12553, A => n12552, ZN => 
                           n12554);
   U6027 : INV_X1 port map( A => n12554, ZN => n12559);
   U6028 : INV_X1 port map( A => n12555, ZN => n12556);
   U6029 : NOR2_X1 port map( A1 => n12557, A2 => n12556, ZN => n12558);
   U6030 : XNOR2_X1 port map( A => n12559, B => n12558, ZN => n8406);
   U6031 : NAND2_X1 port map( A1 => n12560, A2 => n12575, ZN => n12561);
   U6032 : NAND2_X1 port map( A1 => n12561, A2 => n12568, ZN => n12562);
   U6033 : AOI21_X1 port map( B1 => n10707, B2 => n12563, A => n12562, ZN => 
                           n12566);
   U6034 : NAND2_X1 port map( A1 => n12598, A2 => n12603, ZN => n12565);
   U6035 : XNOR2_X1 port map( A => n12566, B => n12565, ZN => I2_dtemp_31_port)
                           ;
   U6036 : INV_X1 port map( A => FP_A(1), ZN => n12567);
   U6037 : XNOR2_X1 port map( A => FP_A(2), B => n12567, ZN => n14701);
   U6038 : NAND2_X1 port map( A1 => n12569, A2 => n12568, ZN => n13774);
   U6039 : NOR2_X1 port map( A1 => n12570, A2 => n13774, ZN => n12572);
   U6040 : AND2_X1 port map( A1 => n13769, A2 => n13767, ZN => n12571);
   U6041 : NAND3_X1 port map( A1 => n13772, A2 => n12572, A3 => n12571, ZN => 
                           n13612);
   U6042 : NAND2_X1 port map( A1 => n12574, A2 => n12573, ZN => n13773);
   U6043 : NOR2_X1 port map( A1 => n13773, A2 => n13774, ZN => n12602);
   U6044 : AND2_X1 port map( A1 => n12577, A2 => n12575, ZN => n12600);
   U6045 : NAND2_X1 port map( A1 => n12600, A2 => n12598, ZN => n13775);
   U6046 : NOR2_X1 port map( A1 => n12602, A2 => n13775, ZN => n12576);
   U6047 : NAND2_X1 port map( A1 => n13612, A2 => n12576, ZN => n13756);
   U6048 : NAND2_X1 port map( A1 => n12585, A2 => n13776, ZN => n12596);
   U6049 : INV_X1 port map( A => n12585, ZN => n12582);
   U6050 : INV_X1 port map( A => n12577, ZN => n12579);
   U6051 : AND2_X1 port map( A1 => n12578, A2 => n12606, ZN => n12604);
   U6052 : OAI21_X1 port map( B1 => n12603, B2 => n12579, A => n12604, ZN => 
                           n13777);
   U6053 : AOI21_X1 port map( B1 => n13777, B2 => n13776, A => n12580, ZN => 
                           n12581);
   U6054 : OAI22_X1 port map( A1 => n13756, A2 => n12596, B1 => n12582, B2 => 
                           n12581, ZN => n12584);
   U6055 : AND2_X1 port map( A1 => n13608, A2 => n12597, ZN => n12583);
   U6056 : XNOR2_X1 port map( A => n12584, B => n12583, ZN => n14937);
   U6057 : NAND2_X1 port map( A1 => n12585, A2 => n12597, ZN => n13764);
   U6058 : NAND3_X1 port map( A1 => n13762, A2 => n13776, A3 => n13758, ZN => 
                           n12586);
   U6059 : NOR2_X1 port map( A1 => n13764, A2 => n12586, ZN => n12589);
   U6060 : INV_X1 port map( A => n12589, ZN => n12592);
   U6061 : NAND2_X1 port map( A1 => n12588, A2 => n12587, ZN => n13792);
   U6062 : AOI21_X1 port map( B1 => n13792, B2 => n13758, A => n13757, ZN => 
                           n12591);
   U6063 : NAND2_X1 port map( A1 => n13777, A2 => n12589, ZN => n12590);
   U6064 : OAI211_X1 port map( C1 => n13756, C2 => n12592, A => n12591, B => 
                           n12590, ZN => n12595);
   U6065 : INV_X1 port map( A => n12423, ZN => n12593);
   U6066 : XNOR2_X1 port map( A => n10817, B => n12593, ZN => n12594);
   U6067 : XNOR2_X1 port map( A => n12595, B => n12594, ZN => I2_dtemp_39_port)
                           ;
   U6068 : NAND2_X1 port map( A1 => n13612, A2 => n12612, ZN => n12615);
   U6069 : INV_X1 port map( A => n12596, ZN => n12599);
   U6070 : NAND4_X1 port map( A1 => n12600, A2 => n12599, A3 => n12598, A4 => 
                           n12597, ZN => n12601);
   U6071 : OR2_X1 port map( A1 => n12602, A2 => n12601, ZN => n13606);
   U6072 : NAND2_X1 port map( A1 => n12604, A2 => n12603, ZN => n12610);
   U6073 : INV_X1 port map( A => n13764, ZN => n12609);
   U6074 : NAND3_X1 port map( A1 => n12607, A2 => n12606, A3 => n12605, ZN => 
                           n12608);
   U6075 : NAND4_X1 port map( A1 => n12610, A2 => n12609, A3 => n13776, A4 => 
                           n12608, ZN => n13609);
   U6076 : NAND2_X1 port map( A1 => n13609, A2 => n12611, ZN => n12613);
   U6077 : NAND2_X1 port map( A1 => n12613, A2 => n12612, ZN => n12614);
   U6078 : OAI21_X1 port map( B1 => n12615, B2 => n13606, A => n12614, ZN => 
                           n12619);
   U6079 : AND2_X1 port map( A1 => n12617, A2 => n12616, ZN => n12618);
   U6080 : XNOR2_X1 port map( A => n12619, B => n12618, ZN => n14933);
   U6081 : NAND2_X1 port map( A1 => n12621, A2 => n12620, ZN => n12624);
   U6082 : INV_X1 port map( A => n12622, ZN => n12623);
   U6083 : OR2_X1 port map( A1 => n10738, A2 => n14447, ZN => n12627);
   U6084 : XNOR2_X1 port map( A => n14593, B => n13277, ZN => n12625);
   U6085 : MUX2_X1 port map( A => n14020, B => n10939, S => n8334, Z => n12629)
                           ;
   U6086 : NAND2_X1 port map( A1 => n14458, A2 => n12230, ZN => n12628);
   U6087 : NAND2_X1 port map( A1 => n12629, A2 => n12628, ZN => n13094);
   U6088 : INV_X1 port map( A => n13094, ZN => n13098);
   U6089 : XNOR2_X1 port map( A => n13097, B => n13098, ZN => n12632);
   U6090 : NAND2_X1 port map( A1 => n12163, A2 => n14719, ZN => n12630);
   U6091 : NAND2_X1 port map( A1 => n12631, A2 => n12630, ZN => n13095);
   U6092 : XNOR2_X1 port map( A => n12632, B => n13095, ZN => n13157);
   U6093 : MUX2_X1 port map( A => n14878, B => n12163, S => n10864, Z => n12634
                           );
   U6094 : MUX2_X1 port map( A => n13915, B => n14779, S => n8329, Z => n12638)
                           ;
   U6095 : XOR2_X1 port map( A => n14720, B => n8325, Z => n12636);
   U6096 : NAND2_X1 port map( A1 => n12636, A2 => n10679, ZN => n12637);
   U6097 : NAND2_X1 port map( A1 => n12638, A2 => n12637, ZN => n13089);
   U6098 : MUX2_X1 port map( A => n10745, B => n12639, S => n14788, Z => n12643
                           );
   U6099 : XNOR2_X1 port map( A => n10905, B => n12671, ZN => n12641);
   U6100 : NAND2_X1 port map( A1 => n12641, A2 => n12640, ZN => n12642);
   U6101 : NAND2_X1 port map( A1 => n12643, A2 => n12642, ZN => n13088);
   U6102 : INV_X1 port map( A => n13158, ZN => n12644);
   U6103 : OAI21_X1 port map( B1 => n13156, B2 => n13157, A => n12644, ZN => 
                           n12646);
   U6104 : NAND2_X1 port map( A1 => n13156, A2 => n13157, ZN => n12645);
   U6105 : AND2_X1 port map( A1 => n12646, A2 => n12645, ZN => n14936);
   U6106 : NOR2_X1 port map( A1 => n13628, A2 => n14596, ZN => n14710);
   U6107 : NAND2_X1 port map( A1 => n14639, A2 => FP_A(19), ZN => n14640);
   U6108 : MUX2_X1 port map( A => n13362, B => n14114, S => n10841, Z => n12647
                           );
   U6109 : INV_X1 port map( A => n12647, ZN => n12649);
   U6110 : MUX2_X1 port map( A => n10713, B => n10636, S => n13261, Z => n12648
                           );
   U6111 : NAND2_X1 port map( A1 => n12649, A2 => n12648, ZN => n12652);
   U6112 : NAND2_X1 port map( A1 => n12652, A2 => n14129, ZN => n12686);
   U6113 : MUX2_X1 port map( A => n14878, B => n11971, S => n14450, Z => n12650
                           );
   U6114 : AND2_X1 port map( A1 => n12651, A2 => n12650, ZN => n14131);
   U6115 : NAND2_X1 port map( A1 => n12686, A2 => n14131, ZN => n12653);
   U6116 : INV_X1 port map( A => n12652, ZN => n14130);
   U6117 : INV_X1 port map( A => n14129, ZN => n12672);
   U6118 : NAND2_X1 port map( A1 => n14130, A2 => n12672, ZN => n12685);
   U6119 : NAND2_X1 port map( A1 => n12653, A2 => n12685, ZN => n12654);
   U6120 : OR2_X1 port map( A1 => intadd_62_SUM_0_port, A2 => n12654, ZN => 
                           n14261);
   U6121 : MUX2_X1 port map( A => n10885, B => n13817, S => n10831, Z => n12656
                           );
   U6122 : MUX2_X1 port map( A => n13819, B => n14882, S => n13234, Z => n12655
                           );
   U6123 : AND2_X1 port map( A1 => n12656, A2 => n12655, ZN => n14161);
   U6124 : INV_X1 port map( A => n14161, ZN => n12660);
   U6125 : MUX2_X1 port map( A => n14114, B => n13362, S => n13261, Z => n12657
                           );
   U6126 : INV_X1 port map( A => n12657, ZN => n12659);
   U6127 : MUX2_X1 port map( A => n10713, B => n10636, S => n13262, Z => n12658
                           );
   U6128 : NAND2_X1 port map( A1 => n12659, A2 => n12658, ZN => n14162);
   U6129 : NAND2_X1 port map( A1 => n12660, A2 => n14162, ZN => n12664);
   U6130 : MUX2_X1 port map( A => n12163, B => n13824, S => n13813, Z => n12661
                           );
   U6131 : NAND2_X1 port map( A1 => n12662, A2 => n12661, ZN => n14163);
   U6132 : INV_X1 port map( A => n14163, ZN => n12663);
   U6133 : NAND2_X1 port map( A1 => n12664, A2 => n12663, ZN => n12667);
   U6134 : INV_X1 port map( A => n14162, ZN => n12665);
   U6135 : NAND2_X1 port map( A1 => n12665, A2 => n14161, ZN => n12666);
   U6136 : NAND2_X1 port map( A1 => n12667, A2 => n12666, ZN => n14159);
   U6137 : INV_X1 port map( A => n14159, ZN => n12683);
   U6138 : MUX2_X1 port map( A => n14840, B => n10645, S => n13450, Z => n12669
                           );
   U6139 : MUX2_X1 port map( A => n10925, B => n10736, S => n10726, Z => n12668
                           );
   U6140 : OAI21_X1 port map( B1 => n14121, B2 => n12669, A => n12668, ZN => 
                           n14150);
   U6141 : INV_X1 port map( A => n14150, ZN => n12670);
   U6142 : INV_X1 port map( A => n12674, ZN => n14149);
   U6143 : NAND2_X1 port map( A1 => n12670, A2 => n14149, ZN => n12678);
   U6144 : NAND3_X1 port map( A1 => n14734, A2 => n14463, A3 => n12671, ZN => 
                           n13000);
   U6145 : NAND2_X1 port map( A1 => n13372, A2 => n13000, ZN => n12673);
   U6146 : MUX2_X1 port map( A => n12673, B => n12672, S => n10841, Z => n14151
                           );
   U6147 : INV_X1 port map( A => n14151, ZN => n12676);
   U6148 : NAND2_X1 port map( A1 => n14150, A2 => n12674, ZN => n12675);
   U6149 : NAND2_X1 port map( A1 => n12676, A2 => n12675, ZN => n12677);
   U6150 : NAND2_X1 port map( A1 => n12678, A2 => n12677, ZN => n14158);
   U6151 : INV_X1 port map( A => n14158, ZN => n12682);
   U6152 : MUX2_X1 port map( A => n14880, B => n10886, S => n13810, Z => n12680
                           );
   U6153 : MUX2_X1 port map( A => n13819, B => n14882, S => n14478, Z => n12679
                           );
   U6154 : AND2_X1 port map( A1 => n12680, A2 => n12679, ZN => n14157);
   U6155 : OAI21_X1 port map( B1 => n14159, B2 => n14158, A => n14157, ZN => 
                           n12681);
   U6156 : OAI21_X1 port map( B1 => n12683, B2 => n12682, A => n12681, ZN => 
                           n14262);
   U6157 : NAND2_X1 port map( A1 => n14261, A2 => n14262, ZN => n12689);
   U6158 : INV_X1 port map( A => n14131, ZN => n12684);
   U6159 : NAND2_X1 port map( A1 => n12685, A2 => n12684, ZN => n12687);
   U6160 : AND2_X1 port map( A1 => n12687, A2 => n12686, ZN => n12688);
   U6161 : NAND2_X1 port map( A1 => intadd_62_SUM_0_port, A2 => n12688, ZN => 
                           n14260);
   U6162 : NAND2_X1 port map( A1 => n12689, A2 => n14260, ZN => n12690);
   U6163 : NAND2_X1 port map( A1 => intadd_62_SUM_1_port, A2 => n12690, ZN => 
                           intadd_61_n6);
   U6164 : NOR2_X1 port map( A1 => intadd_62_SUM_1_port, A2 => n12690, ZN => 
                           intadd_61_n5);
   U6165 : INV_X1 port map( A => intadd_61_n5, ZN => n12691);
   U6166 : NAND2_X1 port map( A1 => n12691, A2 => intadd_61_n6, ZN => 
                           intadd_61_n2);
   U6167 : XNOR2_X1 port map( A => n14708, B => FP_A(7), ZN => n14571);
   U6168 : XNOR2_X1 port map( A => FP_A(13), B => n14661, ZN => n14670);
   U6169 : OR2_X1 port map( A1 => n12692, A2 => n14641, ZN => FP_Z(30));
   U6170 : MUX2_X1 port map( A => n14840, B => n10645, S => n8329, Z => n12694)
                           ;
   U6171 : MUX2_X1 port map( A => n13442, B => n10736, S => n14482, Z => n12693
                           );
   U6172 : OAI21_X1 port map( B1 => n14121, B2 => n12694, A => n12693, ZN => 
                           n12719);
   U6173 : AND2_X1 port map( A1 => n10914, A2 => n13809, ZN => n14142);
   U6174 : XNOR2_X1 port map( A => n12719, B => n14142, ZN => n12696);
   U6175 : NAND2_X1 port map( A1 => n13346, A2 => n14716, ZN => n12695);
   U6176 : MUX2_X1 port map( A => n12695, B => n14134, S => n10841, Z => n12716
                           );
   U6177 : XNOR2_X1 port map( A => n12696, B => n12716, ZN => n12712);
   U6178 : MUX2_X1 port map( A => n13372, B => n13371, S => n13262, Z => n12698
                           );
   U6179 : MUX2_X1 port map( A => n12142, B => n10641, S => n13823, Z => n12697
                           );
   U6180 : NAND2_X1 port map( A1 => n12698, A2 => n12697, ZN => n12760);
   U6181 : MUX2_X1 port map( A => n13817, B => n10885, S => n10742, Z => n12700
                           );
   U6182 : MUX2_X1 port map( A => n13819, B => n14882, S => n10913, Z => n12699
                           );
   U6183 : NAND2_X1 port map( A1 => n12700, A2 => n12699, ZN => n12759);
   U6184 : INV_X1 port map( A => n12759, ZN => n12701);
   U6185 : NAND2_X1 port map( A1 => n13449, A2 => n14492, ZN => n12758);
   U6186 : NAND2_X1 port map( A1 => n12701, A2 => n12758, ZN => n12704);
   U6187 : INV_X1 port map( A => n12758, ZN => n12702);
   U6188 : AND2_X1 port map( A1 => n12759, A2 => n12702, ZN => n12703);
   U6189 : AOI21_X1 port map( B1 => n12760, B2 => n12704, A => n12703, ZN => 
                           n12713);
   U6190 : NAND2_X1 port map( A1 => n12712, A2 => n12713, ZN => n14225);
   U6191 : MUX2_X1 port map( A => n14114, B => n13362, S => n13823, Z => n12706
                           );
   U6192 : MUX2_X1 port map( A => n12146, B => n11225, S => n10631, Z => n12705
                           );
   U6193 : NOR2_X1 port map( A1 => n12706, A2 => n12705, ZN => n12832);
   U6194 : MUX2_X1 port map( A => n13372, B => n13371, S => n13261, Z => n12708
                           );
   U6195 : MUX2_X1 port map( A => n13000, B => n12142, S => n14467, Z => n12707
                           );
   U6196 : AND2_X1 port map( A1 => n12708, A2 => n12707, ZN => n12831);
   U6197 : MUX2_X1 port map( A => n12163, B => n14878, S => n13234, Z => n12709
                           );
   U6198 : AND2_X1 port map( A1 => n12710, A2 => n12709, ZN => n12830);
   U6199 : INV_X1 port map( A => n14226, ZN => n12711);
   U6200 : NAND2_X1 port map( A1 => n14225, A2 => n12711, ZN => n12727);
   U6201 : INV_X1 port map( A => n12712, ZN => n12715);
   U6202 : INV_X1 port map( A => n12713, ZN => n12714);
   U6203 : NAND2_X1 port map( A1 => n12715, A2 => n12714, ZN => n14224);
   U6204 : INV_X1 port map( A => n12716, ZN => n12718);
   U6205 : INV_X1 port map( A => n14142, ZN => n14140);
   U6206 : NAND2_X1 port map( A1 => n12719, A2 => n14140, ZN => n12717);
   U6207 : NAND2_X1 port map( A1 => n12718, A2 => n12717, ZN => n14169);
   U6208 : INV_X1 port map( A => n12719, ZN => n12720);
   U6209 : NAND2_X1 port map( A1 => n12720, A2 => n14142, ZN => n14168);
   U6210 : NAND2_X1 port map( A1 => n14169, A2 => n14168, ZN => n12726);
   U6211 : MUX2_X1 port map( A => n13824, B => n12163, S => n10831, Z => n12721
                           );
   U6212 : NAND2_X1 port map( A1 => n12722, A2 => n12721, ZN => n14171);
   U6213 : MUX2_X1 port map( A => n14880, B => n10886, S => n13234, Z => n12724
                           );
   U6214 : MUX2_X1 port map( A => n13819, B => n14882, S => n14449, Z => n12723
                           );
   U6215 : NAND2_X1 port map( A1 => n12724, A2 => n12723, ZN => n14170);
   U6216 : XNOR2_X1 port map( A => n14171, B => n14170, ZN => n12725);
   U6217 : XNOR2_X1 port map( A => n12726, B => n12725, ZN => n12728);
   U6218 : NAND3_X1 port map( A1 => n12727, A2 => n14224, A3 => n12728, ZN => 
                           n14235);
   U6219 : NAND2_X1 port map( A1 => n14224, A2 => n14226, ZN => n12730);
   U6220 : INV_X1 port map( A => n12728, ZN => n12729);
   U6221 : NAND3_X1 port map( A1 => n12730, A2 => n12729, A3 => n14225, ZN => 
                           n14234);
   U6222 : NAND2_X1 port map( A1 => n14235, A2 => n14234, ZN => n12749);
   U6223 : MUX2_X1 port map( A => n14114, B => n13362, S => n8325, Z => n12731)
                           ;
   U6224 : INV_X1 port map( A => n12731, ZN => n12733);
   U6225 : MUX2_X1 port map( A => n10713, B => n10636, S => n8329, Z => n12732)
                           ;
   U6226 : NAND2_X1 port map( A1 => n12733, A2 => n12732, ZN => n12755);
   U6227 : MUX2_X1 port map( A => n14840, B => n10645, S => n13813, Z => n12735
                           );
   U6228 : MUX2_X1 port map( A => n10925, B => n10738, S => n10831, Z => n12734
                           );
   U6229 : OAI21_X1 port map( B1 => n14121, B2 => n12735, A => n12734, ZN => 
                           n12754);
   U6230 : NAND2_X1 port map( A1 => n12755, A2 => n12754, ZN => n12739);
   U6231 : MUX2_X1 port map( A => n13824, B => n12163, S => n14945, Z => n12736
                           );
   U6232 : NAND2_X1 port map( A1 => n12737, A2 => n12736, ZN => n12756);
   U6233 : INV_X1 port map( A => n12756, ZN => n12738);
   U6234 : NAND2_X1 port map( A1 => n12739, A2 => n12738, ZN => n12740);
   U6235 : OAI21_X1 port map( B1 => n12755, B2 => n12754, A => n12740, ZN => 
                           n12751);
   U6236 : MUX2_X1 port map( A => n10885, B => n13817, S => n14945, Z => n12742
                           );
   U6237 : MUX2_X1 port map( A => n13819, B => n14882, S => n10743, Z => n12741
                           );
   U6238 : AND2_X1 port map( A1 => n12742, A2 => n12741, ZN => n12750);
   U6239 : MUX2_X1 port map( A => n12805, B => n13346, S => n10841, Z => n12795
                           );
   U6240 : MUX2_X1 port map( A => n13283, B => n14716, S => n13261, Z => n12794
                           );
   U6241 : NAND2_X1 port map( A1 => n12795, A2 => n12794, ZN => n12746);
   U6242 : AND2_X1 port map( A1 => n13328, A2 => n13809, ZN => n12801);
   U6243 : INV_X1 port map( A => n12801, ZN => n12803);
   U6244 : NAND2_X1 port map( A1 => n12743, A2 => n13809, ZN => n12744);
   U6245 : NAND2_X1 port map( A1 => n12803, A2 => n12744, ZN => n12791);
   U6246 : OR2_X1 port map( A1 => n12803, A2 => n14457, ZN => n12792);
   U6247 : INV_X1 port map( A => n12792, ZN => n12745);
   U6248 : AOI21_X1 port map( B1 => n12746, B2 => n12791, A => n12745, ZN => 
                           n12752);
   U6249 : OAI21_X1 port map( B1 => n12751, B2 => n12750, A => n12752, ZN => 
                           n12748);
   U6250 : NAND2_X1 port map( A1 => n12751, A2 => n12750, ZN => n12747);
   U6251 : AND2_X1 port map( A1 => n12748, A2 => n12747, ZN => n14232);
   U6252 : XNOR2_X1 port map( A => n12749, B => n14232, ZN => n14870);
   U6253 : INV_X1 port map( A => n14870, ZN => n14871);
   U6254 : XNOR2_X1 port map( A => n12751, B => n12750, ZN => n12753);
   U6255 : XNOR2_X1 port map( A => n12753, B => n12752, ZN => n12814);
   U6256 : INV_X1 port map( A => n12814, ZN => n12779);
   U6257 : XNOR2_X1 port map( A => n12755, B => n12754, ZN => n12757);
   U6258 : XNOR2_X1 port map( A => n12757, B => n12756, ZN => n13309);
   U6259 : XNOR2_X1 port map( A => n12759, B => n12758, ZN => n12761);
   U6260 : XNOR2_X1 port map( A => n12761, B => n12760, ZN => n13307);
   U6261 : INV_X1 port map( A => n13307, ZN => n12775);
   U6262 : MUX2_X1 port map( A => n13346, B => n12805, S => n13262, Z => n12763
                           );
   U6263 : MUX2_X1 port map( A => n13347, B => n14716, S => n13823, Z => n12762
                           );
   U6264 : NAND2_X1 port map( A1 => n12763, A2 => n12762, ZN => n13382);
   U6265 : AND2_X1 port map( A1 => n13368, A2 => B_SIG_8_port, ZN => n13379);
   U6266 : OAI21_X1 port map( B1 => n12764, B2 => n11703, A => n13809, ZN => 
                           n13380);
   U6267 : INV_X1 port map( A => n13380, ZN => n12765);
   U6268 : OAI21_X1 port map( B1 => n13382, B2 => n13379, A => n12765, ZN => 
                           n13300);
   U6269 : MUX2_X1 port map( A => n13372, B => n13371, S => n13823, Z => n12767
                           );
   U6270 : MUX2_X1 port map( A => n10745, B => n13373, S => n10726, Z => n12766
                           );
   U6271 : NAND2_X1 port map( A1 => n12767, A2 => n12766, ZN => n13299);
   U6272 : INV_X1 port map( A => n13299, ZN => n12768);
   U6273 : NAND2_X1 port map( A1 => n13300, A2 => n12768, ZN => n12771);
   U6274 : MUX2_X1 port map( A => n13817, B => n10885, S => n10913, Z => n12770
                           );
   U6275 : MUX2_X1 port map( A => n13819, B => n14882, S => n13327, Z => n12769
                           );
   U6276 : NAND2_X1 port map( A1 => n12770, A2 => n12769, ZN => n13298);
   U6277 : NAND2_X1 port map( A1 => n12771, A2 => n13298, ZN => n12774);
   U6278 : INV_X1 port map( A => n13300, ZN => n12772);
   U6279 : NAND2_X1 port map( A1 => n12772, A2 => n13299, ZN => n12773);
   U6280 : NAND2_X1 port map( A1 => n12774, A2 => n12773, ZN => n13308);
   U6281 : OAI21_X1 port map( B1 => n13309, B2 => n12775, A => n13308, ZN => 
                           n12777);
   U6282 : NAND2_X1 port map( A1 => n13309, A2 => n12775, ZN => n12776);
   U6283 : NAND2_X1 port map( A1 => n12779, A2 => n12778, ZN => n14228);
   U6284 : MUX2_X1 port map( A => n14114, B => n13362, S => n8329, Z => n12780)
                           ;
   U6285 : INV_X1 port map( A => n12780, ZN => n12782);
   U6286 : MUX2_X1 port map( A => n10713, B => n10636, S => n13239, Z => n12781
                           );
   U6287 : MUX2_X1 port map( A => n14878, B => n12163, S => n14477, Z => n12785
                           );
   U6288 : NAND2_X1 port map( A1 => n12786, A2 => n12785, ZN => n13296);
   U6289 : INV_X1 port map( A => n13296, ZN => n12787);
   U6290 : NAND2_X1 port map( A1 => n12788, A2 => n13294, ZN => n12789);
   U6291 : NAND2_X1 port map( A1 => n12790, A2 => n12789, ZN => n13254);
   U6292 : INV_X1 port map( A => n13254, ZN => n12798);
   U6293 : NAND2_X1 port map( A1 => n12792, A2 => n12791, ZN => n12793);
   U6294 : AND3_X1 port map( A1 => n12795, A2 => n12794, A3 => n12793, ZN => 
                           n12797);
   U6295 : AOI21_X1 port map( B1 => n12795, B2 => n12794, A => n12793, ZN => 
                           n12796);
   U6296 : NAND2_X1 port map( A1 => n12798, A2 => n13255, ZN => n12812);
   U6297 : MUX2_X1 port map( A => n10645, B => n14840, S => n10831, Z => n12800
                           );
   U6298 : MUX2_X1 port map( A => n10925, B => n10736, S => n14452, Z => n12799
                           );
   U6299 : OAI21_X1 port map( B1 => n14121, B2 => n12800, A => n12799, ZN => 
                           n12804);
   U6300 : INV_X1 port map( A => n12804, ZN => n12802);
   U6301 : NAND2_X1 port map( A1 => n12802, A2 => n12801, ZN => n13226);
   U6302 : NAND2_X1 port map( A1 => n12804, A2 => n12803, ZN => n13225);
   U6303 : MUX2_X1 port map( A => n13346, B => n11651, S => n13261, Z => n12807
                           );
   U6304 : MUX2_X1 port map( A => n13283, B => n14716, S => n8334, Z => n12806)
                           ;
   U6305 : NAND2_X1 port map( A1 => n13225, A2 => n12808, ZN => n12809);
   U6306 : NAND2_X1 port map( A1 => n13226, A2 => n12809, ZN => n13253);
   U6307 : INV_X1 port map( A => n13255, ZN => n12811);
   U6308 : AOI22_X1 port map( A1 => n12812, A2 => n13253, B1 => n12811, B2 => 
                           n13254, ZN => n14230);
   U6309 : INV_X1 port map( A => n14230, ZN => n12813);
   U6310 : NAND2_X1 port map( A1 => n14228, A2 => n12813, ZN => n12816);
   U6311 : NAND2_X1 port map( A1 => n12815, A2 => n12814, ZN => n14229);
   U6312 : NAND2_X1 port map( A1 => n12816, A2 => n14229, ZN => n14252);
   U6313 : MUX2_X1 port map( A => n14114, B => n13362, S => n13262, Z => n12817
                           );
   U6314 : INV_X1 port map( A => n12817, ZN => n12819);
   U6315 : MUX2_X1 port map( A => n10713, B => n10636, S => n13823, Z => n12818
                           );
   U6316 : NAND2_X1 port map( A1 => n12819, A2 => n12818, ZN => n14135);
   U6317 : XNOR2_X1 port map( A => n14135, B => n14134, ZN => n12822);
   U6318 : MUX2_X1 port map( A => n13371, B => n13372, S => n10841, Z => n12821
                           );
   U6319 : MUX2_X1 port map( A => n13373, B => n13000, S => n13261, Z => n12820
                           );
   U6320 : NAND2_X1 port map( A1 => n12821, A2 => n12820, ZN => n14137);
   U6321 : XNOR2_X1 port map( A => n12822, B => n14137, ZN => n12826);
   U6322 : MUX2_X1 port map( A => n14840, B => n10645, S => n10631, Z => n12824
                           );
   U6323 : MUX2_X1 port map( A => n13442, B => n10736, S => n14450, Z => n12823
                           );
   U6324 : OAI21_X1 port map( B1 => n14121, B2 => n12824, A => n12823, ZN => 
                           n14143);
   U6325 : AND2_X1 port map( A1 => n10742, A2 => n10702, ZN => n14144);
   U6326 : XNOR2_X1 port map( A => n14144, B => n14140, ZN => n12825);
   U6327 : XNOR2_X1 port map( A => n14143, B => n12825, ZN => n12827);
   U6328 : NAND2_X1 port map( A1 => n12826, A2 => n12827, ZN => n14238);
   U6329 : INV_X1 port map( A => n12826, ZN => n12829);
   U6330 : INV_X1 port map( A => n12827, ZN => n12828);
   U6331 : NAND2_X1 port map( A1 => n12829, A2 => n12828, ZN => n14177);
   U6332 : NAND2_X1 port map( A1 => n14238, A2 => n14177, ZN => n12833);
   U6333 : FA_X1 port map( A => n12832, B => n12831, CI => n12830, CO => n14176
                           , S => n14226);
   U6334 : XNOR2_X1 port map( A => n12833, B => n14176, ZN => n14251);
   U6335 : NAND2_X1 port map( A1 => n14252, A2 => n14251, ZN => n14873);
   U6336 : NAND2_X1 port map( A1 => n14873, A2 => n14870, ZN => n14852);
   U6337 : NAND2_X1 port map( A1 => FP_A(3), A2 => FP_A(4), ZN => n14699);
   U6338 : NOR2_X1 port map( A1 => n12835, A2 => n12834, ZN => n12836);
   U6339 : NOR2_X1 port map( A1 => intadd_58_A_1_port, A2 => n12836, ZN => 
                           n13903);
   U6340 : MUX2_X1 port map( A => n13979, B => n13908, S => n8401, Z => n12840)
                           ;
   U6341 : MUX2_X1 port map( A => n13920, B => n14728, S => n14465, Z => n12838
                           );
   U6342 : INV_X1 port map( A => n12838, ZN => n12839);
   U6343 : OR2_X1 port map( A1 => n12840, A2 => n12839, ZN => n12967);
   U6344 : MUX2_X1 port map( A => n10680, B => n11043, S => n14025, Z => n12842
                           );
   U6345 : MUX2_X1 port map( A => n10725, B => n11834, S => n14777, Z => n12841
                           );
   U6346 : NAND2_X1 port map( A1 => n12842, A2 => n12841, ZN => n13940);
   U6347 : MUX2_X1 port map( A => n14020, B => n10940, S => B_SIG_8_port, Z => 
                           n12844);
   U6348 : NAND2_X1 port map( A1 => n14451, A2 => n14771, ZN => n12843);
   U6349 : NAND2_X1 port map( A1 => n12844, A2 => n12843, ZN => n13938);
   U6350 : INV_X1 port map( A => n13938, ZN => n12845);
   U6351 : NAND2_X1 port map( A1 => n14813, A2 => n14719, ZN => n13937);
   U6352 : NAND2_X1 port map( A1 => n12845, A2 => n13937, ZN => n12846);
   U6353 : NAND2_X1 port map( A1 => n13940, A2 => n12846, ZN => n12849);
   U6354 : INV_X1 port map( A => n13937, ZN => n12847);
   U6355 : NAND2_X1 port map( A1 => n12847, A2 => n13938, ZN => n12848);
   U6356 : NAND2_X1 port map( A1 => n12849, A2 => n12848, ZN => n12966);
   U6357 : OAI21_X1 port map( B1 => n13903, B2 => n12967, A => n12966, ZN => 
                           n12851);
   U6358 : NAND2_X1 port map( A1 => n13903, A2 => n12967, ZN => n12850);
   U6359 : NAND2_X1 port map( A1 => n12851, A2 => n12850, ZN => n12983);
   U6360 : MUX2_X1 port map( A => n13979, B => n13908, S => n13924, Z => n12854
                           );
   U6361 : MUX2_X1 port map( A => n13920, B => n14728, S => n14448, Z => n12852
                           );
   U6362 : INV_X1 port map( A => n12852, ZN => n12853);
   U6363 : MUX2_X1 port map( A => n14017, B => n11201, S => B_SIG_8_port, Z => 
                           n12856);
   U6364 : MUX2_X1 port map( A => n13915, B => n14779, S => n13485, Z => n12855
                           );
   U6365 : AND2_X1 port map( A1 => n12856, A2 => n12855, ZN => n12868);
   U6366 : INV_X1 port map( A => n12868, ZN => n12857);
   U6367 : XNOR2_X1 port map( A => n12870, B => n12857, ZN => n12861);
   U6368 : MUX2_X1 port map( A => n13323, B => n11743, S => n14025, Z => n12858
                           );
   U6369 : INV_X1 port map( A => n12858, ZN => n12860);
   U6370 : MUX2_X1 port map( A => n10640, B => n13868, S => n14594, Z => n12859
                           );
   U6371 : NAND2_X1 port map( A1 => n12860, A2 => n12859, ZN => n12871);
   U6372 : XNOR2_X1 port map( A => n12861, B => n12871, ZN => n12982);
   U6373 : FA_X1 port map( A => n12983, B => n12982, CI => intadd_58_SUM_1_port
                           , CO => n12986, S => n_1343);
   U6374 : XNOR2_X1 port map( A => n12862, B => n13174, ZN => n12863);
   U6375 : XNOR2_X1 port map( A => n12863, B => n13173, ZN => n13168);
   U6376 : NAND2_X1 port map( A1 => n12865, A2 => n12864, ZN => n12867);
   U6377 : XNOR2_X1 port map( A => n12867, B => n12866, ZN => n13170);
   U6378 : INV_X1 port map( A => n13170, ZN => n12891);
   U6379 : NAND2_X1 port map( A1 => n12870, A2 => n12871, ZN => n12869);
   U6380 : NAND2_X1 port map( A1 => n12869, A2 => n12868, ZN => n12875);
   U6381 : INV_X1 port map( A => n12870, ZN => n12873);
   U6382 : INV_X1 port map( A => n12871, ZN => n12872);
   U6383 : NAND2_X1 port map( A1 => n12873, A2 => n12872, ZN => n12874);
   U6384 : NAND2_X1 port map( A1 => n12875, A2 => n12874, ZN => n13856);
   U6385 : NAND2_X1 port map( A1 => n12877, A2 => n12876, ZN => n12879);
   U6386 : XNOR2_X1 port map( A => n12879, B => n12878, ZN => n12888);
   U6387 : MUX2_X1 port map( A => n11043, B => n11957, S => n8350, Z => n12881)
                           ;
   U6388 : MUX2_X1 port map( A => n10725, B => n11834, S => n14785, Z => n12880
                           );
   U6389 : AND2_X1 port map( A1 => n12881, A2 => n12880, ZN => n13864);
   U6390 : MUX2_X1 port map( A => n14020, B => n10939, S => n8351, Z => n12883)
                           ;
   U6391 : NAND2_X1 port map( A1 => n14453, A2 => n14771, ZN => n12882);
   U6392 : NAND2_X1 port map( A1 => n12883, A2 => n12882, ZN => n13861);
   U6393 : AND2_X1 port map( A1 => n14727, A2 => n14719, ZN => n12884);
   U6394 : NAND2_X1 port map( A1 => n13861, A2 => n12884, ZN => n12886);
   U6395 : INV_X1 port map( A => n13861, ZN => n12885);
   U6396 : INV_X1 port map( A => n12884, ZN => n13862);
   U6397 : AOI22_X1 port map( A1 => n13864, A2 => n12886, B1 => n12885, B2 => 
                           n13862, ZN => n12887);
   U6398 : NAND2_X1 port map( A1 => n12888, A2 => n12887, ZN => n13857);
   U6399 : NAND2_X1 port map( A1 => n13856, A2 => n13857, ZN => n12890);
   U6400 : INV_X1 port map( A => n12887, ZN => n12889);
   U6401 : NAND2_X1 port map( A1 => n12889, A2 => n10715, ZN => n13858);
   U6402 : NAND2_X1 port map( A1 => n12890, A2 => n13858, ZN => n13169);
   U6403 : XNOR2_X1 port map( A => n12891, B => n13169, ZN => n12892);
   U6404 : XNOR2_X1 port map( A => n13168, B => n12892, ZN => n13617);
   U6405 : OAI22_X1 port map( A1 => intadd_58_SUM_2_port, A2 => n12986, B1 => 
                           intadd_58_n1, B2 => n13617, ZN => n12893);
   U6406 : INV_X1 port map( A => n12893, ZN => n14745);
   U6407 : NAND2_X1 port map( A1 => n12894, A2 => n12895, ZN => n12896);
   U6408 : INV_X1 port map( A => n12894, ZN => n12904);
   U6409 : INV_X1 port map( A => n12895, ZN => n12905);
   U6410 : AOI22_X1 port map( A1 => n12906, A2 => n12896, B1 => n12904, B2 => 
                           n12905, ZN => n12903);
   U6411 : AOI21_X1 port map( B1 => n12898, B2 => n12897, A => n12900, ZN => 
                           n12899);
   U6412 : INV_X1 port map( A => n12899, ZN => n12902);
   U6413 : OR2_X1 port map( A1 => n12903, A2 => n12909, ZN => n13121);
   U6414 : OAI21_X1 port map( B1 => n12906, B2 => n12905, A => n12904, ZN => 
                           n12908);
   U6415 : NAND2_X1 port map( A1 => n12906, A2 => n12905, ZN => n12907);
   U6416 : NAND2_X1 port map( A1 => n12940, A2 => n12910, ZN => n12912);
   U6417 : NAND2_X1 port map( A1 => n12912, A2 => n12911, ZN => n13123);
   U6418 : NAND2_X1 port map( A1 => n13121, A2 => n12913, ZN => n12920);
   U6419 : XNOR2_X1 port map( A => n12914, B => n12915, ZN => n12919);
   U6420 : AND2_X1 port map( A1 => n12917, A2 => n12916, ZN => n12918);
   U6421 : XNOR2_X1 port map( A => n12919, B => n12918, ZN => n13127);
   U6422 : XNOR2_X1 port map( A => n12920, B => n13127, ZN => n12952);
   U6423 : INV_X1 port map( A => n13128, ZN => n12925);
   U6424 : XNOR2_X1 port map( A => n12952, B => n12925, ZN => n12930);
   U6425 : NAND2_X1 port map( A1 => n12927, A2 => n12926, ZN => n12929);
   U6426 : XNOR2_X1 port map( A => n12929, B => n12928, ZN => n12953);
   U6427 : NAND2_X1 port map( A1 => n12930, A2 => n12953, ZN => n13575);
   U6428 : INV_X1 port map( A => n13123, ZN => n12931);
   U6429 : XNOR2_X1 port map( A => n12932, B => n12931, ZN => n12948);
   U6430 : NAND2_X1 port map( A1 => n12934, A2 => n12933, ZN => n12937);
   U6432 : NAND2_X1 port map( A1 => n12937, A2 => n12935, ZN => n12947);
   U6433 : NAND2_X1 port map( A1 => n12948, A2 => n12947, ZN => n14068);
   U6434 : XNOR2_X1 port map( A => n12939, B => n12938, ZN => n12944);
   U6435 : XNOR2_X1 port map( A => n12941, B => n12940, ZN => n12943);
   U6436 : OAI21_X1 port map( B1 => n12944, B2 => n12943, A => n12942, ZN => 
                           n12946);
   U6437 : NAND2_X1 port map( A1 => n12944, A2 => n12943, ZN => n12945);
   U6438 : NAND2_X1 port map( A1 => n12946, A2 => n12945, ZN => n14070);
   U6439 : NAND2_X1 port map( A1 => n14068, A2 => n14070, ZN => n12951);
   U6440 : INV_X1 port map( A => n12947, ZN => n12950);
   U6441 : INV_X1 port map( A => n12948, ZN => n12949);
   U6442 : NAND2_X1 port map( A1 => n12950, A2 => n12949, ZN => n14069);
   U6443 : NAND2_X1 port map( A1 => n12951, A2 => n14069, ZN => n13577);
   U6444 : NAND2_X1 port map( A1 => n13575, A2 => n13577, ZN => n12956);
   U6445 : XNOR2_X1 port map( A => n10916, B => n12952, ZN => n12955);
   U6446 : INV_X1 port map( A => n12953, ZN => n12954);
   U6447 : NAND2_X1 port map( A1 => n12955, A2 => n12954, ZN => n13576);
   U6448 : NAND2_X1 port map( A1 => n12956, A2 => n13576, ZN => n14803);
   U6449 : XNOR2_X1 port map( A => n12958, B => n12957, ZN => n12959);
   U6450 : XNOR2_X1 port map( A => n12959, B => n12960, ZN => n12989);
   U6451 : NAND2_X1 port map( A1 => n12962, A2 => n12961, ZN => n12965);
   U6452 : INV_X1 port map( A => n12963, ZN => n12964);
   U6453 : XNOR2_X1 port map( A => n12965, B => n12964, ZN => n12988);
   U6454 : OR2_X1 port map( A1 => n12989, A2 => n12988, ZN => n14764);
   U6455 : XNOR2_X1 port map( A => n12967, B => n12966, ZN => n13901);
   U6456 : XNOR2_X1 port map( A => n13901, B => n13903, ZN => n12980);
   U6457 : OR2_X1 port map( A1 => intadd_58_SUM_0_port, A2 => n12980, ZN => 
                           n12981);
   U6458 : MUX2_X1 port map( A => n13979, B => n13908, S => n13914, Z => n12970
                           );
   U6459 : MUX2_X1 port map( A => n13920, B => n14728, S => n14593, Z => n12968
                           );
   U6460 : INV_X1 port map( A => n12968, ZN => n12969);
   U6461 : OR2_X1 port map( A1 => n12970, A2 => n12969, ZN => n13936);
   U6462 : MUX2_X1 port map( A => n10680, B => n11043, S => n14594, Z => n12972
                           );
   U6463 : MUX2_X1 port map( A => n10725, B => n11834, S => n14719, Z => n12971
                           );
   U6464 : NAND2_X1 port map( A1 => n12972, A2 => n12971, ZN => n13918);
   U6465 : OAI21_X1 port map( B1 => n11043, B2 => n14719, A => n10725, ZN => 
                           n13919);
   U6466 : NAND2_X1 port map( A1 => n13918, A2 => n13919, ZN => n13947);
   U6467 : MUX2_X1 port map( A => n14017, B => n13984, S => n13924, Z => n12974
                           );
   U6468 : MUX2_X1 port map( A => n13915, B => n14779, S => n14731, Z => n12973
                           );
   U6469 : AND2_X1 port map( A1 => n12974, A2 => n12973, ZN => n12976);
   U6470 : NAND2_X1 port map( A1 => n13947, A2 => n12976, ZN => n12975);
   U6471 : NAND2_X1 port map( A1 => n13936, A2 => n12975, ZN => n12979);
   U6472 : INV_X1 port map( A => n13947, ZN => n12977);
   U6473 : INV_X1 port map( A => n12976, ZN => n13935);
   U6474 : NAND2_X1 port map( A1 => n12977, A2 => n13935, ZN => n12978);
   U6475 : NAND2_X1 port map( A1 => n12979, A2 => n12978, ZN => n13904);
   U6476 : AOI22_X1 port map( A1 => n12981, A2 => n13904, B1 => n12980, B2 => 
                           intadd_58_SUM_0_port, ZN => n14058);
   U6477 : INV_X1 port map( A => n12982, ZN => n12984);
   U6478 : XNOR2_X1 port map( A => n12984, B => n12983, ZN => n12985);
   U6479 : XNOR2_X1 port map( A => intadd_58_SUM_1_port, B => n12985, ZN => 
                           n14059);
   U6480 : NAND2_X1 port map( A1 => intadd_58_SUM_2_port, A2 => n12986, ZN => 
                           n12987);
   U6481 : OAI21_X1 port map( B1 => n14058, B2 => n14059, A => n12987, ZN => 
                           n14747);
   U6482 : NAND2_X1 port map( A1 => n12989, A2 => n12988, ZN => n13167);
   U6483 : NAND2_X1 port map( A1 => n13167, A2 => n12990, ZN => n14763);
   U6484 : XNOR2_X1 port map( A => n12994, B => n12993, ZN => n13559);
   U6486 : XNOR2_X1 port map( A => n12997, B => n12996, ZN => n12999);
   U6487 : XNOR2_X1 port map( A => n12999, B => n12998, ZN => n14081);
   U6488 : NAND2_X1 port map( A1 => n14079, A2 => n14081, ZN => n13034);
   U6489 : INV_X1 port map( A => n13000, ZN => n13001);
   U6490 : AOI22_X1 port map( A1 => n10637, A2 => n14464, B1 => n13001, B2 => 
                           n8351, ZN => n13003);
   U6491 : NAND2_X1 port map( A1 => n13003, A2 => n13002, ZN => n13004);
   U6492 : NAND2_X1 port map( A1 => n13004, A2 => n13005, ZN => n13009);
   U6493 : INV_X1 port map( A => n13005, ZN => n13008);
   U6494 : XNOR2_X1 port map( A => n13010, B => n11594, ZN => n13011);
   U6495 : XNOR2_X1 port map( A => n13012, B => n13011, ZN => n13136);
   U6496 : INV_X1 port map( A => n13136, ZN => n13023);
   U6497 : NAND2_X1 port map( A1 => n13016, A2 => n13017, ZN => n13015);
   U6498 : NAND2_X1 port map( A1 => n13015, A2 => n13014, ZN => n13021);
   U6499 : INV_X1 port map( A => n13016, ZN => n13019);
   U6500 : INV_X1 port map( A => n13017, ZN => n13018);
   U6501 : NAND2_X1 port map( A1 => n13019, A2 => n13018, ZN => n13020);
   U6502 : NAND2_X1 port map( A1 => n13021, A2 => n13020, ZN => n13137);
   U6503 : INV_X1 port map( A => n13137, ZN => n13022);
   U6504 : OAI21_X1 port map( B1 => n13138, B2 => n13023, A => n13022, ZN => 
                           n13025);
   U6505 : NAND2_X1 port map( A1 => n13138, A2 => n13023, ZN => n13024);
   U6506 : NAND2_X1 port map( A1 => n13025, A2 => n13024, ZN => n14078);
   U6507 : INV_X1 port map( A => n14078, ZN => n13033);
   U6508 : INV_X1 port map( A => n14081, ZN => n13032);
   U6509 : INV_X1 port map( A => n13026, ZN => n13027);
   U6510 : NAND2_X1 port map( A1 => n13028, A2 => n13027, ZN => n13029);
   U6511 : AND2_X1 port map( A1 => n10694, A2 => n13029, ZN => n13031);
   U6512 : AND2_X1 port map( A1 => n13558, A2 => n13559, ZN => n14200);
   U6513 : XNOR2_X1 port map( A => n13036, B => n10698, ZN => n13148);
   U6514 : XNOR2_X1 port map( A => n13037, B => n13038, ZN => n13039);
   U6515 : XNOR2_X1 port map( A => n13039, B => n13040, ZN => n13147);
   U6516 : XNOR2_X1 port map( A => n13042, B => n13041, ZN => n13044);
   U6517 : XNOR2_X1 port map( A => n13044, B => n13043, ZN => n13146);
   U6518 : INV_X1 port map( A => n13146, ZN => n13045);
   U6519 : OAI21_X1 port map( B1 => n13148, B2 => n13147, A => n13045, ZN => 
                           n13047);
   U6520 : NAND2_X1 port map( A1 => n13148, A2 => n13147, ZN => n13046);
   U6521 : NAND2_X1 port map( A1 => n13047, A2 => n13046, ZN => n14202);
   U6522 : XNOR2_X1 port map( A => n13048, B => n13049, ZN => n13053);
   U6523 : XNOR2_X1 port map( A => n13051, B => n13050, ZN => n13052);
   U6524 : XNOR2_X1 port map( A => n13053, B => n13052, ZN => n13550);
   U6525 : INV_X1 port map( A => n13550, ZN => n14201);
   U6526 : XNOR2_X1 port map( A => n13056, B => n13055, ZN => n13565);
   U6527 : NAND2_X1 port map( A1 => n13058, A2 => n13057, ZN => n13060);
   U6528 : XNOR2_X1 port map( A => n13060, B => n13059, ZN => n13564);
   U6529 : XNOR2_X1 port map( A => n13564, B => n13565, ZN => n13065);
   U6530 : XNOR2_X1 port map( A => n13062, B => n13061, ZN => n13064);
   U6531 : XNOR2_X1 port map( A => n13064, B => n13063, ZN => n13566);
   U6532 : INV_X1 port map( A => n13558, ZN => n13066);
   U6533 : NAND2_X1 port map( A1 => n10947, A2 => n13066, ZN => n14206);
   U6534 : OAI21_X1 port map( B1 => n13560, B2 => n14200, A => n14206, ZN => 
                           n14827);
   U6535 : XNOR2_X1 port map( A => n13067, B => n13068, ZN => n13070);
   U6536 : XNOR2_X1 port map( A => n13070, B => n13069, ZN => n13557);
   U6537 : INV_X1 port map( A => n13557, ZN => n13083);
   U6538 : OAI21_X1 port map( B1 => n13072, B2 => n13073, A => n13071, ZN => 
                           n13075);
   U6539 : NAND2_X1 port map( A1 => n13073, A2 => n13072, ZN => n13074);
   U6540 : NAND2_X1 port map( A1 => n13075, A2 => n13074, ZN => n13554);
   U6541 : INV_X1 port map( A => n13554, ZN => n13082);
   U6542 : NAND2_X1 port map( A1 => n13077, A2 => n13076, ZN => n13079);
   U6543 : XNOR2_X1 port map( A => n13079, B => n13078, ZN => n13555);
   U6544 : NAND2_X1 port map( A1 => n13557, A2 => n13555, ZN => n13081);
   U6545 : NAND2_X1 port map( A1 => n13555, A2 => n13554, ZN => n13080);
   U6546 : OAI211_X1 port map( C1 => n13083, C2 => n13082, A => n13081, B => 
                           n13080, ZN => n13129);
   U6547 : XNOR2_X1 port map( A => n13085, B => n13084, ZN => n13087);
   U6548 : XNOR2_X1 port map( A => n13087, B => n13086, ZN => n13130);
   U6549 : OR2_X1 port map( A1 => n13129, A2 => n13130, ZN => n14073);
   U6550 : NAND2_X1 port map( A1 => n13089, A2 => n13088, ZN => n13090);
   U6551 : AND2_X1 port map( A1 => n13093, A2 => n13092, ZN => n13102);
   U6552 : NAND2_X1 port map( A1 => n13097, A2 => n13094, ZN => n13096);
   U6553 : NAND2_X1 port map( A1 => n13096, A2 => n13095, ZN => n13101);
   U6554 : INV_X1 port map( A => n13097, ZN => n13099);
   U6555 : NAND2_X1 port map( A1 => n13099, A2 => n13098, ZN => n13100);
   U6556 : NAND2_X1 port map( A1 => n13101, A2 => n13100, ZN => n13154);
   U6557 : NAND2_X1 port map( A1 => n13152, A2 => n13154, ZN => n13105);
   U6558 : INV_X1 port map( A => n13102, ZN => n13103);
   U6559 : NAND2_X1 port map( A1 => n13104, A2 => n13103, ZN => n13153);
   U6560 : NAND2_X1 port map( A1 => n13105, A2 => n13153, ZN => n13193);
   U6561 : XNOR2_X1 port map( A => n13107, B => n13106, ZN => n13116);
   U6562 : XNOR2_X1 port map( A => n13116, B => n13115, ZN => n13114);
   U6563 : XNOR2_X1 port map( A => n13109, B => n13108, ZN => n13113);
   U6564 : XNOR2_X1 port map( A => n10915, B => n13110, ZN => n13112);
   U6565 : XNOR2_X1 port map( A => n13113, B => n13112, ZN => n13117);
   U6566 : NAND2_X1 port map( A1 => n13114, A2 => n13117, ZN => n13191);
   U6567 : NAND2_X1 port map( A1 => n13193, A2 => n13191, ZN => n13120);
   U6568 : XOR2_X1 port map( A => n13116, B => n13115, Z => n13119);
   U6569 : INV_X1 port map( A => n13117, ZN => n13118);
   U6570 : NAND2_X1 port map( A1 => n13119, A2 => n13118, ZN => n13192);
   U6571 : NAND2_X1 port map( A1 => n13120, A2 => n13192, ZN => n14075);
   U6572 : NAND2_X1 port map( A1 => n14073, A2 => n14075, ZN => n13151);
   U6573 : NAND2_X1 port map( A1 => n13128, A2 => n13127, ZN => n13124);
   U6574 : INV_X1 port map( A => n13121, ZN => n13122);
   U6575 : NAND2_X1 port map( A1 => n13124, A2 => n13122, ZN => n13126);
   U6576 : INV_X1 port map( A => n13215, ZN => n13131);
   U6577 : NAND2_X1 port map( A1 => n13129, A2 => n13130, ZN => n14074);
   U6578 : INV_X1 port map( A => n13216, ZN => n14098);
   U6579 : XNOR2_X1 port map( A => n13137, B => n13136, ZN => n13139);
   U6580 : XNOR2_X1 port map( A => n13139, B => n13138, ZN => n14189);
   U6581 : NAND2_X1 port map( A1 => n13140, A2 => n13141, ZN => n13145);
   U6582 : INV_X1 port map( A => n13141, ZN => n13142);
   U6583 : XNOR2_X1 port map( A => n14189, B => n14188, ZN => n13150);
   U6584 : XNOR2_X1 port map( A => n13147, B => n13146, ZN => n13149);
   U6585 : XNOR2_X1 port map( A => n13149, B => n13148, ZN => n14190);
   U6586 : XNOR2_X1 port map( A => n13150, B => n10918, ZN => n14097);
   U6587 : NAND2_X1 port map( A1 => n13151, A2 => n14074, ZN => n13217);
   U6588 : NAND2_X1 port map( A1 => n13217, A2 => n13215, ZN => n14099);
   U6589 : OAI211_X1 port map( C1 => n14100, C2 => n14098, A => n14097, B => 
                           n14099, ZN => n14793);
   U6590 : AND2_X1 port map( A1 => n13153, A2 => n13152, ZN => n13155);
   U6591 : XOR2_X1 port map( A => n13155, B => n13154, Z => intadd_46_A_2_port)
                           ;
   U6592 : INV_X1 port map( A => n14755, ZN => n14756);
   U6593 : XNOR2_X1 port map( A => n13157, B => n13158, ZN => n13159);
   U6594 : XNOR2_X1 port map( A => n13159, B => n13156, ZN => n14066);
   U6595 : NAND2_X1 port map( A1 => intadd_46_SUM_1_port, A2 => n14066, ZN => 
                           n13164);
   U6596 : NAND2_X1 port map( A1 => n13164, A2 => n13163, ZN => n13166);
   U6597 : OR2_X1 port map( A1 => intadd_46_SUM_1_port, A2 => n14066, ZN => 
                           n13165);
   U6598 : NAND2_X1 port map( A1 => n13166, A2 => n13165, ZN => n14796);
   U6599 : XNOR2_X1 port map( A => n10820, B => n10765, ZN => n14772);
   U6600 : NAND2_X1 port map( A1 => n13167, A2 => n14764, ZN => n14766);
   U6601 : FA_X1 port map( A => n13170, B => n13169, CI => n13168, CO => n13602
                           , S => n_1344);
   U6602 : INV_X1 port map( A => n13171, ZN => n13178);
   U6605 : XNOR2_X1 port map( A => n13177, B => n13178, ZN => n13601);
   U6606 : NAND2_X1 port map( A1 => n13602, A2 => n13601, ZN => n14751);
   U6607 : NAND2_X1 port map( A1 => n13180, A2 => n13179, ZN => n13182);
   U6608 : XNOR2_X1 port map( A => n13182, B => n13181, ZN => 
                           intadd_58_A_2_port);
   U6609 : XNOR2_X1 port map( A => n13183, B => n13184, ZN => n13185);
   U6610 : XNOR2_X1 port map( A => n13185, B => n13186, ZN => 
                           intadd_66_B_1_port);
   U6611 : NAND2_X1 port map( A1 => n10919, A2 => n13220, ZN => n13190);
   U6612 : XNOR2_X1 port map( A => n13190, B => n13219, ZN => n13528);
   U6613 : INV_X1 port map( A => n13528, ZN => n14802);
   U6614 : NAND2_X1 port map( A1 => n13192, A2 => n13191, ZN => n13194);
   U6615 : XNOR2_X1 port map( A => n13194, B => n13193, ZN => 
                           intadd_46_A_3_port);
   U6616 : INV_X1 port map( A => n13195, ZN => n13198);
   U6617 : XNOR2_X1 port map( A => intadd_56_A_3_port, B => n13196, ZN => 
                           n13197);
   U6618 : XNOR2_X1 port map( A => n13198, B => n13197, ZN => n14758);
   U6619 : INV_X1 port map( A => n13199, ZN => n13205);
   U6620 : INV_X1 port map( A => n13200, ZN => n13201);
   U6621 : NOR2_X1 port map( A1 => n13205, A2 => n13201, ZN => n13203);
   U6622 : NAND2_X1 port map( A1 => n13203, A2 => n13202, ZN => n13208);
   U6623 : INV_X1 port map( A => n13204, ZN => n13207);
   U6624 : AOI22_X1 port map( A1 => n13208, A2 => n13207, B1 => n13206, B2 => 
                           n13205, ZN => intadd_46_B_1_port);
   U6625 : XNOR2_X1 port map( A => n10740, B => n13210, ZN => n13211);
   U6626 : XNOR2_X1 port map( A => n13211, B => n13212, ZN => n14829);
   U6627 : INV_X1 port map( A => n14827, ZN => n13213);
   U6628 : NAND2_X1 port map( A1 => n13213, A2 => n14829, ZN => n14828);
   U6629 : INV_X1 port map( A => n13214, ZN => n14794);
   U6630 : NAND2_X1 port map( A1 => n10820, A2 => n10813, ZN => n14776);
   U6631 : XNOR2_X1 port map( A => n13216, B => n13215, ZN => n13218);
   U6632 : XNOR2_X1 port map( A => n10839, B => n10838, ZN => n14804);
   U6633 : OAI21_X1 port map( B1 => n14100, B2 => n14098, A => n14099, ZN => 
                           n14810);
   U6634 : NAND2_X1 port map( A1 => n10919, A2 => n13219, ZN => n13222);
   U6635 : AOI21_X1 port map( B1 => n13222, B2 => n13220, A => n14092, ZN => 
                           n13224);
   U6636 : INV_X1 port map( A => n14092, ZN => n13223);
   U6637 : OAI22_X1 port map( A1 => n13224, A2 => n13551, B1 => n13223, B2 => 
                           n10727, ZN => n14807);
   U6638 : NAND2_X1 port map( A1 => n13226, A2 => n13225, ZN => n13227);
   U6639 : INV_X1 port map( A => n13394, ZN => n13252);
   U6640 : MUX2_X1 port map( A => n14878, B => n12163, S => n14455, Z => n13245
                           );
   U6641 : NAND2_X1 port map( A1 => n13246, A2 => n13245, ZN => n13231);
   U6642 : INV_X1 port map( A => n13228, ZN => n13229);
   U6643 : OR2_X1 port map( A1 => n11743, A2 => n13229, ZN => n13244);
   U6644 : INV_X1 port map( A => n13244, ZN => n13230);
   U6645 : NAND2_X1 port map( A1 => n13231, A2 => n13230, ZN => n13317);
   U6646 : MUX2_X1 port map( A => n13448, B => n13449, S => n10841, Z => n13233
                           );
   U6647 : MUX2_X1 port map( A => n14833, B => n13451, S => n13261, Z => n13232
                           );
   U6648 : AND2_X1 port map( A1 => n13233, A2 => n13232, ZN => n13319);
   U6649 : NAND2_X1 port map( A1 => n13317, A2 => n13319, ZN => n13248);
   U6650 : MUX2_X1 port map( A => n14840, B => n10645, S => n13234, Z => n13236
                           );
   U6651 : MUX2_X1 port map( A => n13442, B => n10736, S => n10869, Z => n13235
                           );
   U6652 : OAI21_X1 port map( B1 => n14121, B2 => n13236, A => n13235, ZN => 
                           n13243);
   U6653 : MUX2_X1 port map( A => n13372, B => n13371, S => n10631, Z => n13238
                           );
   U6654 : MUX2_X1 port map( A => n10641, B => n12142, S => n14450, Z => n13237
                           );
   U6655 : NAND2_X1 port map( A1 => n13238, A2 => n13237, ZN => n13242);
   U6656 : INV_X1 port map( A => n13406, ZN => n13383);
   U6657 : MUX2_X1 port map( A => n14114, B => n13362, S => n13239, Z => n13241
                           );
   U6658 : MUX2_X1 port map( A => n12146, B => n11225, S => n14478, Z => n13240
                           );
   U6659 : NOR2_X1 port map( A1 => n13241, A2 => n13240, ZN => n13403);
   U6660 : NAND2_X1 port map( A1 => n13383, A2 => n13403, ZN => n13247);
   U6661 : NOR2_X1 port map( A1 => n13243, A2 => n13242, ZN => n13404);
   U6662 : INV_X1 port map( A => n13404, ZN => n13384);
   U6663 : NAND3_X1 port map( A1 => n13246, A2 => n13245, A3 => n13244, ZN => 
                           n13318);
   U6664 : NAND4_X1 port map( A1 => n13248, A2 => n13247, A3 => n13384, A4 => 
                           n13318, ZN => n13389);
   U6665 : INV_X1 port map( A => n13403, ZN => n13385);
   U6666 : NAND2_X1 port map( A1 => n10692, A2 => n13385, ZN => n13407);
   U6667 : INV_X1 port map( A => n13319, ZN => n13249);
   U6668 : NAND2_X1 port map( A1 => n13318, A2 => n13249, ZN => n13250);
   U6669 : NAND4_X1 port map( A1 => n13407, A2 => n13250, A3 => n13317, A4 => 
                           n13383, ZN => n13390);
   U6670 : INV_X1 port map( A => n13390, ZN => n13251);
   U6671 : AOI21_X1 port map( B1 => n13252, B2 => n13389, A => n13251, ZN => 
                           n13257);
   U6672 : XNOR2_X1 port map( A => n13253, B => n13254, ZN => n13256);
   U6673 : XNOR2_X1 port map( A => n13256, B => n13255, ZN => n13258);
   U6674 : NAND2_X1 port map( A1 => n13257, A2 => n13258, ZN => n14221);
   U6675 : INV_X1 port map( A => n13389, ZN => n13259);
   U6676 : AOI21_X1 port map( B1 => n13394, B2 => n13390, A => n13259, ZN => 
                           n13260);
   U6677 : NAND2_X1 port map( A1 => n10912, A2 => n13260, ZN => n14222);
   U6678 : NAND2_X1 port map( A1 => n14221, A2 => n14222, ZN => n13306);
   U6679 : MUX2_X1 port map( A => n13449, B => n13448, S => n13261, Z => n13264
                           );
   U6680 : MUX2_X1 port map( A => n14833, B => n12783, S => n13262, Z => n13263
                           );
   U6681 : NAND2_X1 port map( A1 => n13264, A2 => n13263, ZN => n13272);
   U6682 : INV_X1 port map( A => n13272, ZN => n13270);
   U6683 : MUX2_X1 port map( A => n10640, B => n13266, S => n10841, Z => n13267
                           );
   U6684 : NAND2_X1 port map( A1 => n13268, A2 => n13267, ZN => n13271);
   U6685 : INV_X1 port map( A => n13271, ZN => n13269);
   U6686 : NAND2_X1 port map( A1 => n13270, A2 => n13269, ZN => n13419);
   U6687 : NAND2_X1 port map( A1 => n13272, A2 => n13271, ZN => n13418);
   U6688 : MUX2_X1 port map( A => n12163, B => n13824, S => n13273, Z => n13274
                           );
   U6689 : AND2_X1 port map( A1 => n13275, A2 => n13274, ZN => n13420);
   U6690 : NAND2_X1 port map( A1 => n13418, A2 => n13420, ZN => n13276);
   U6691 : NAND2_X1 port map( A1 => n13419, A2 => n13276, ZN => n13315);
   U6692 : MUX2_X1 port map( A => n10925, B => n10738, S => n14477, Z => n13281
                           );
   U6693 : XNOR2_X1 port map( A => n13277, B => n10869, ZN => n13278);
   U6694 : NAND2_X1 port map( A1 => n13279, A2 => n13278, ZN => n13280);
   U6695 : NAND2_X1 port map( A1 => n13281, A2 => n13280, ZN => n13413);
   U6696 : MUX2_X1 port map( A => n13283, B => n14716, S => n13282, Z => n13286
                           );
   U6697 : XNOR2_X1 port map( A => n13823, B => n10877, ZN => n13284);
   U6698 : NAND2_X1 port map( A1 => n13285, A2 => n13286, ZN => n13412);
   U6699 : NAND2_X1 port map( A1 => B_SIG_8_port, A2 => n13809, ZN => n13411);
   U6700 : AOI21_X1 port map( B1 => n13412, B2 => n13413, A => n13411, ZN => 
                           n13288);
   U6701 : NOR2_X1 port map( A1 => n10719, A2 => n13413, ZN => n13287);
   U6702 : NOR2_X1 port map( A1 => n13288, A2 => n13287, ZN => n13292);
   U6703 : MUX2_X1 port map( A => n14880, B => n10885, S => n13327, Z => n13290
                           );
   U6704 : MUX2_X1 port map( A => n13819, B => n14882, S => n13328, Z => n13289
                           );
   U6705 : NAND2_X1 port map( A1 => n13290, A2 => n13289, ZN => n13291);
   U6706 : NAND2_X1 port map( A1 => n13292, A2 => n13291, ZN => n13314);
   U6707 : INV_X1 port map( A => n13313, ZN => n13293);
   U6708 : AOI21_X1 port map( B1 => n13315, B2 => n13314, A => n13293, ZN => 
                           n13727);
   U6709 : XNOR2_X1 port map( A => n13295, B => n13294, ZN => n13297);
   U6710 : XNOR2_X1 port map( A => n13297, B => n13296, ZN => n13304);
   U6711 : INV_X1 port map( A => n13304, ZN => n13301);
   U6712 : NAND2_X1 port map( A1 => n13301, A2 => n10710, ZN => n13724);
   U6713 : INV_X1 port map( A => n13724, ZN => n13302);
   U6714 : NAND2_X1 port map( A1 => n13304, A2 => n13303, ZN => n13725);
   U6715 : NAND2_X1 port map( A1 => n13305, A2 => n13725, ZN => n14220);
   U6716 : XNOR2_X1 port map( A => n13306, B => n14220, ZN => n13312);
   U6717 : XNOR2_X1 port map( A => n13307, B => n13308, ZN => n13310);
   U6718 : XNOR2_X1 port map( A => n13310, B => n13309, ZN => n13311);
   U6719 : NAND2_X1 port map( A1 => n10734, A2 => n13311, ZN => n14845);
   U6720 : NAND2_X1 port map( A1 => n10769, A2 => n10829, ZN => n14842);
   U6721 : NAND2_X1 port map( A1 => n13314, A2 => n13313, ZN => n13316);
   U6722 : XNOR2_X1 port map( A => n13316, B => n13315, ZN => n13360);
   U6723 : INV_X1 port map( A => n13360, ZN => n13322);
   U6724 : NAND2_X1 port map( A1 => n13318, A2 => n13317, ZN => n13320);
   U6725 : XNOR2_X1 port map( A => n13320, B => n13319, ZN => n13359);
   U6726 : INV_X1 port map( A => n13359, ZN => n13321);
   U6727 : NAND2_X1 port map( A1 => n13322, A2 => n13321, ZN => n14215);
   U6728 : MUX2_X1 port map( A => n11743, B => n13323, S => n14726, Z => n13324
                           );
   U6729 : INV_X1 port map( A => n13324, ZN => n13326);
   U6730 : MUX2_X1 port map( A => n10640, B => n13868, S => n14459, Z => n13325
                           );
   U6731 : NAND2_X1 port map( A1 => n13326, A2 => n13325, ZN => n13531);
   U6732 : MUX2_X1 port map( A => n12163, B => n13824, S => n13328, Z => n13329
                           );
   U6733 : NAND2_X1 port map( A1 => n13330, A2 => n13329, ZN => n13530);
   U6734 : NAND2_X1 port map( A1 => n13531, A2 => n13530, ZN => n13337);
   U6735 : MUX2_X1 port map( A => n14114, B => n13362, S => n13234, Z => n13331
                           );
   U6736 : INV_X1 port map( A => n13331, ZN => n13333);
   U6737 : MUX2_X1 port map( A => n10713, B => n10636, S => n14449, Z => n13332
                           );
   U6738 : NAND2_X1 port map( A1 => n13333, A2 => n13332, ZN => n13529);
   U6739 : INV_X1 port map( A => n13529, ZN => n13336);
   U6740 : INV_X1 port map( A => n13531, ZN => n13335);
   U6741 : INV_X1 port map( A => n13530, ZN => n13334);
   U6742 : AOI22_X1 port map( A1 => n13337, A2 => n13336, B1 => n13335, B2 => 
                           n13334, ZN => n13345);
   U6743 : MUX2_X1 port map( A => n14840, B => n10645, S => n10742, Z => n13338
                           );
   U6744 : INV_X1 port map( A => n13338, ZN => n13339);
   U6745 : NAND2_X1 port map( A1 => n13339, A2 => n14460, ZN => n13341);
   U6746 : MUX2_X1 port map( A => n10925, B => n10738, S => n14455, Z => n13340
                           );
   U6747 : NAND2_X1 port map( A1 => n13341, A2 => n13340, ZN => n13424);
   U6748 : NAND2_X1 port map( A1 => n13924, A2 => n13809, ZN => n13643);
   U6749 : INV_X1 port map( A => n13643, ZN => n13458);
   U6750 : NAND2_X1 port map( A1 => n13424, A2 => n13458, ZN => n13343);
   U6751 : NAND2_X1 port map( A1 => n10905, A2 => n14718, ZN => n13422);
   U6752 : AND2_X1 port map( A1 => n13340, A2 => n13643, ZN => n13342);
   U6753 : AOI22_X1 port map( A1 => n13343, A2 => n13422, B1 => n13342, B2 => 
                           n13341, ZN => n13344);
   U6754 : OR2_X1 port map( A1 => n13345, A2 => n13344, ZN => n13464);
   U6755 : NAND2_X1 port map( A1 => n13345, A2 => n13344, ZN => n13465);
   U6756 : MUX2_X1 port map( A => n13346, B => n12805, S => n10631, Z => n13349
                           );
   U6757 : MUX2_X1 port map( A => n13347, B => n14716, S => n11649, Z => n13348
                           );
   U6758 : NAND2_X1 port map( A1 => n13349, A2 => n13348, ZN => n13535);
   U6759 : INV_X1 port map( A => n13535, ZN => n13353);
   U6760 : MUX2_X1 port map( A => n13372, B => n13371, S => n13810, Z => n13351
                           );
   U6761 : MUX2_X1 port map( A => n10745, B => n12142, S => n10831, Z => n13350
                           );
   U6762 : AND2_X1 port map( A1 => n13351, A2 => n13350, ZN => n13355);
   U6763 : INV_X1 port map( A => n13355, ZN => n13352);
   U6764 : NAND2_X1 port map( A1 => n14507, A2 => n8355, ZN => n13516);
   U6765 : NAND2_X1 port map( A1 => n13352, A2 => n13516, ZN => n13533);
   U6766 : NAND2_X1 port map( A1 => n13353, A2 => n13533, ZN => n13356);
   U6767 : INV_X1 port map( A => n13516, ZN => n13354);
   U6768 : NAND2_X1 port map( A1 => n13355, A2 => n13354, ZN => n13534);
   U6769 : NAND2_X1 port map( A1 => n13356, A2 => n13534, ZN => n13466);
   U6770 : NAND2_X1 port map( A1 => n13465, A2 => n13466, ZN => n13357);
   U6771 : AND2_X1 port map( A1 => n13464, A2 => n13357, ZN => n14217);
   U6772 : INV_X1 port map( A => n14217, ZN => n13358);
   U6773 : NAND2_X1 port map( A1 => n14215, A2 => n13358, ZN => n13361);
   U6774 : NAND2_X1 port map( A1 => n13360, A2 => n13359, ZN => n14216);
   U6775 : NAND2_X1 port map( A1 => n13361, A2 => n14216, ZN => n13401);
   U6776 : MUX2_X1 port map( A => n13362, B => n14114, S => n10831, Z => n13363
                           );
   U6777 : INV_X1 port map( A => n13363, ZN => n13366);
   U6778 : MUX2_X1 port map( A => n10713, B => n10636, S => n13364, Z => n13365
                           );
   U6779 : NAND2_X1 port map( A1 => n13366, A2 => n13365, ZN => n13417);
   U6780 : MUX2_X1 port map( A => n13817, B => n10885, S => n8351, Z => n13370)
                           ;
   U6781 : MUX2_X1 port map( A => n13819, B => n14882, S => n13368, Z => n13369
                           );
   U6782 : NAND2_X1 port map( A1 => n13370, A2 => n13369, ZN => n13415);
   U6783 : NAND2_X1 port map( A1 => n13417, A2 => n13415, ZN => n13378);
   U6784 : MUX2_X1 port map( A => n13372, B => n13371, S => n8329, Z => n13375)
                           ;
   U6785 : MUX2_X1 port map( A => n13373, B => n10745, S => n13813, Z => n13374
                           );
   U6786 : AND2_X1 port map( A1 => n13375, A2 => n13374, ZN => n13416);
   U6787 : INV_X1 port map( A => n13417, ZN => n13377);
   U6788 : INV_X1 port map( A => n13415, ZN => n13376);
   U6789 : NOR2_X1 port map( A1 => n13380, A2 => n13379, ZN => n13381);
   U6790 : XNOR2_X1 port map( A => n13382, B => n13381, ZN => n13409);
   U6791 : INV_X1 port map( A => n13409, ZN => n13388);
   U6792 : NAND2_X1 port map( A1 => n13384, A2 => n13383, ZN => n13386);
   U6793 : XNOR2_X1 port map( A => n13386, B => n13385, ZN => n13387);
   U6794 : NAND2_X1 port map( A1 => n13390, A2 => n13389, ZN => n13393);
   U6795 : XNOR2_X1 port map( A => n13394, B => n13393, ZN => n13391);
   U6796 : NAND2_X1 port map( A1 => n13392, A2 => n13391, ZN => n13400);
   U6797 : NAND2_X1 port map( A1 => n13401, A2 => n13400, ZN => n13397);
   U6798 : INV_X1 port map( A => n13392, ZN => n13396);
   U6799 : XOR2_X1 port map( A => n13394, B => n13393, Z => n13395);
   U6800 : NAND2_X1 port map( A1 => n13396, A2 => n13395, ZN => n13399);
   U6801 : NAND2_X1 port map( A1 => n13397, A2 => n13399, ZN => n14844);
   U6802 : NAND2_X1 port map( A1 => n13398, A2 => n14844, ZN => n14846);
   U6803 : NAND2_X1 port map( A1 => n13400, A2 => n13399, ZN => n13402);
   U6804 : XNOR2_X1 port map( A => n13402, B => n13401, ZN => n14839);
   U6805 : OAI21_X1 port map( B1 => n13404, B2 => n13406, A => n13403, ZN => 
                           n13405);
   U6806 : OAI21_X1 port map( B1 => n13407, B2 => n13406, A => n13405, ZN => 
                           n13408);
   U6807 : XNOR2_X1 port map( A => n13410, B => n13409, ZN => n13719);
   U6808 : INV_X1 port map( A => n13413, ZN => n13414);
   U6809 : NAND2_X1 port map( A1 => n13419, A2 => n13418, ZN => n13421);
   U6810 : XNOR2_X1 port map( A => n13421, B => n13420, ZN => n13668);
   U6811 : XNOR2_X1 port map( A => n13719, B => n13721, ZN => n13478);
   U6812 : XNOR2_X1 port map( A => n13422, B => n13458, ZN => n13423);
   U6813 : XNOR2_X1 port map( A => n13424, B => n13423, ZN => n13634);
   U6814 : NAND2_X1 port map( A1 => n13426, A2 => n13630, ZN => n13425);
   U6815 : INV_X1 port map( A => n13629, ZN => n13631);
   U6816 : NAND2_X1 port map( A1 => n13425, A2 => n13631, ZN => n13428);
   U6817 : INV_X1 port map( A => n13630, ZN => n13632);
   U6818 : NAND2_X1 port map( A1 => n10703, A2 => n13632, ZN => n13427);
   U6819 : NAND2_X1 port map( A1 => n13428, A2 => n13427, ZN => n13438);
   U6820 : INV_X1 port map( A => n13433, ZN => n13434);
   U6821 : NAND2_X1 port map( A1 => n13634, A2 => n13438, ZN => n13439);
   U6822 : MUX2_X1 port map( A => n14840, B => n10645, S => n10913, Z => n13444
                           );
   U6823 : MUX2_X1 port map( A => n10925, B => n10736, S => n14457, Z => n13443
                           );
   U6824 : NAND2_X1 port map( A1 => n14717, A2 => n14597, ZN => n13445);
   U6825 : MUX2_X1 port map( A => n11834, B => n13445, S => n10841, Z => n13447
                           );
   U6826 : NAND2_X1 port map( A1 => n13447, A2 => n11043, ZN => n13644);
   U6827 : NOR2_X1 port map( A1 => n13651, A2 => n13644, ZN => n13460);
   U6828 : MUX2_X1 port map( A => n13449, B => n13448, S => n13262, Z => n13453
                           );
   U6829 : MUX2_X1 port map( A => n14833, B => n13451, S => n13450, Z => n13452
                           );
   U6830 : NAND2_X1 port map( A1 => n13453, A2 => n13452, ZN => n13656);
   U6831 : INV_X1 port map( A => n13656, ZN => n13454);
   U6832 : NAND2_X1 port map( A1 => n13651, A2 => n13644, ZN => n13459);
   U6833 : OAI211_X1 port map( C1 => n13460, C2 => n13458, A => n13454, B => 
                           n13459, ZN => n13469);
   U6834 : MUX2_X1 port map( A => n14880, B => n10885, S => n12764, Z => n13457
                           );
   U6835 : MUX2_X1 port map( A => n13819, B => n14882, S => B_SIG_8_port, Z => 
                           n13456);
   U6836 : NAND2_X1 port map( A1 => n13457, A2 => n13456, ZN => n13650);
   U6837 : NAND2_X1 port map( A1 => n13469, A2 => n13650, ZN => n13463);
   U6838 : NAND2_X1 port map( A1 => n13459, A2 => n13458, ZN => n13462);
   U6839 : INV_X1 port map( A => n13460, ZN => n13461);
   U6840 : NAND3_X1 port map( A1 => n13462, A2 => n13461, A3 => n13656, ZN => 
                           n13468);
   U6841 : NAND2_X1 port map( A1 => n13463, A2 => n13468, ZN => n13676);
   U6842 : NAND2_X1 port map( A1 => n13677, A2 => n13676, ZN => n13473);
   U6843 : NAND2_X1 port map( A1 => n13465, A2 => n13464, ZN => n13467);
   U6844 : XNOR2_X1 port map( A => n13467, B => n13466, ZN => n13678);
   U6845 : NAND2_X1 port map( A1 => n13473, A2 => n13678, ZN => n13472);
   U6846 : INV_X1 port map( A => n13677, ZN => n13675);
   U6847 : INV_X1 port map( A => n13650, ZN => n13647);
   U6848 : NAND2_X1 port map( A1 => n13468, A2 => n13647, ZN => n13470);
   U6849 : AND2_X1 port map( A1 => n13470, A2 => n13469, ZN => n13674);
   U6850 : INV_X1 port map( A => n13674, ZN => n13474);
   U6851 : NAND2_X1 port map( A1 => n13675, A2 => n13474, ZN => n13471);
   U6852 : NAND2_X1 port map( A1 => n13472, A2 => n13471, ZN => n13723);
   U6853 : AND2_X1 port map( A1 => n13678, A2 => n13473, ZN => n13476);
   U6854 : AND2_X1 port map( A1 => n13675, A2 => n13474, ZN => n13475);
   U6855 : OAI21_X1 port map( B1 => n13476, B2 => n13475, A => n13478, ZN => 
                           n13477);
   U6856 : OAI21_X1 port map( B1 => n13478, B2 => n13723, A => n13477, ZN => 
                           n14850);
   U6857 : NAND2_X1 port map( A1 => n8401, A2 => n8350, ZN => n13479);
   U6858 : NAND3_X1 port map( A1 => n13481, A2 => n13480, A3 => n13479, ZN => 
                           n13484);
   U6859 : AOI21_X1 port map( B1 => n14448, B2 => n14465, A => n13482, ZN => 
                           n13483);
   U6860 : NAND2_X1 port map( A1 => n13484, A2 => n13483, ZN => n13492);
   U6861 : INV_X1 port map( A => n13492, ZN => n13490);
   U6862 : MUX2_X1 port map( A => n14487, B => n13367, S => B_SIG_8_port, Z => 
                           n13488);
   U6863 : MUX2_X1 port map( A => n13486, B => n14480, S => n10904, Z => n13487
                           );
   U6864 : NOR2_X1 port map( A1 => n13488, A2 => n13487, ZN => n13491);
   U6865 : INV_X1 port map( A => n13491, ZN => n13489);
   U6866 : NAND2_X1 port map( A1 => n13490, A2 => n13489, ZN => n13540);
   U6867 : NAND2_X1 port map( A1 => n13492, A2 => n13491, ZN => n13542);
   U6868 : NAND2_X1 port map( A1 => n13540, A2 => n13542, ZN => n13498);
   U6870 : NAND2_X1 port map( A1 => n13495, A2 => n10603, ZN => n13496);
   U6871 : XNOR2_X1 port map( A => n13498, B => n13539, ZN => n13597);
   U6872 : INV_X1 port map( A => n13597, ZN => n13520);
   U6873 : OAI21_X1 port map( B1 => n10924, B2 => n13501, A => n13500, ZN => 
                           n13503);
   U6874 : NAND2_X1 port map( A1 => n10924, A2 => n13501, ZN => n13502);
   U6875 : NAND2_X1 port map( A1 => n13503, A2 => n13502, ZN => n13598);
   U6876 : AND2_X1 port map( A1 => n13505, A2 => n13506, ZN => n13508);
   U6877 : INV_X1 port map( A => n13509, ZN => n13514);
   U6878 : NAND2_X1 port map( A1 => n13510, A2 => n13968, ZN => n13513);
   U6879 : INV_X1 port map( A => n13510, ZN => n13512);
   U6880 : INV_X1 port map( A => n13968, ZN => n13511);
   U6881 : XNOR2_X1 port map( A => n13651, B => n13643, ZN => n13518);
   U6882 : NOR2_X1 port map( A1 => n10638, A2 => n10642, ZN => n13515);
   U6883 : MUX2_X1 port map( A => n13516, B => n13515, S => n14881, Z => n13517
                           );
   U6884 : XNOR2_X1 port map( A => n13518, B => n13517, ZN => n13637);
   U6885 : NAND2_X1 port map( A1 => n13522, A2 => n13521, ZN => n13524);
   U6886 : NAND2_X1 port map( A1 => n13524, A2 => n13523, ZN => n13546);
   U6887 : XNOR2_X1 port map( A => n13549, B => n13546, ZN => n14859);
   U6888 : NOR2_X1 port map( A1 => n13618, A2 => n13601, ZN => n13526);
   U6889 : NOR2_X1 port map( A1 => n10849, A2 => n10848, ZN => n14744);
   U6890 : XNOR2_X1 port map( A => n10764, B => n10867, ZN => n14805);
   U6891 : XNOR2_X1 port map( A => n13530, B => n13529, ZN => n13532);
   U6892 : XNOR2_X1 port map( A => n13531, B => n13532, ZN => n13538);
   U6893 : NAND2_X1 port map( A1 => n13534, A2 => n13533, ZN => n13536);
   U6894 : XNOR2_X1 port map( A => n13536, B => n13535, ZN => n13537);
   U6895 : NAND2_X1 port map( A1 => n13538, A2 => n13537, ZN => n13665);
   U6896 : OR2_X1 port map( A1 => n13538, A2 => n13537, ZN => n13666);
   U6897 : NAND2_X1 port map( A1 => n13665, A2 => n13666, ZN => n13544);
   U6898 : AND2_X1 port map( A1 => n13543, A2 => n13542, ZN => n13663);
   U6899 : XNOR2_X1 port map( A => n13544, B => n13663, ZN => n14858);
   U6900 : INV_X1 port map( A => n13546, ZN => n13545);
   U6901 : NOR2_X1 port map( A1 => n14858, A2 => n13545, ZN => n13548);
   U6902 : INV_X1 port map( A => n14858, ZN => n13547);
   U6903 : OAI22_X1 port map( A1 => n13549, A2 => n13548, B1 => n13547, B2 => 
                           n13546, ZN => n14868);
   U6904 : NAND2_X1 port map( A1 => FP_A(15), A2 => FP_A(16), ZN => n14601);
   U6905 : INV_X1 port map( A => n14094, ZN => n13553);
   U6906 : XNOR2_X1 port map( A => n13550, B => n14202, ZN => n14185);
   U6907 : XNOR2_X1 port map( A => n14185, B => n14207, ZN => n14095);
   U6908 : INV_X1 port map( A => n14095, ZN => n13552);
   U6909 : NAND2_X1 port map( A1 => n14811, A2 => n13551, ZN => n14093);
   U6910 : OAI211_X1 port map( C1 => n13553, C2 => n14092, A => n13552, B => 
                           n14093, ZN => n14791);
   U6911 : XNOR2_X1 port map( A => n13555, B => n13554, ZN => n13556);
   U6912 : XNOR2_X1 port map( A => n13557, B => n13556, ZN => 
                           intadd_46_B_3_port);
   U6913 : XNOR2_X1 port map( A => n13559, B => n13558, ZN => n13561);
   U6914 : XNOR2_X1 port map( A => n13561, B => n13560, ZN => n13574);
   U6915 : OAI21_X1 port map( B1 => n13566, B2 => n13565, A => n13564, ZN => 
                           n13568);
   U6916 : NAND2_X1 port map( A1 => n13566, A2 => n13565, ZN => n13567);
   U6917 : NAND2_X1 port map( A1 => n13568, A2 => n13567, ZN => n13580);
   U6918 : NAND2_X1 port map( A1 => n13569, A2 => n13570, ZN => n13572);
   U6919 : XNOR2_X1 port map( A => n13572, B => n13571, ZN => n13581);
   U6920 : XNOR2_X1 port map( A => n13580, B => n13581, ZN => n13573);
   U6921 : XNOR2_X1 port map( A => n13579, B => n13573, ZN => n14187);
   U6922 : NAND2_X1 port map( A1 => n10859, A2 => n10858, ZN => n14823);
   U6923 : INV_X1 port map( A => n13574, ZN => n14815);
   U6924 : NAND2_X1 port map( A1 => n13576, A2 => n13575, ZN => n13578);
   U6926 : NAND2_X1 port map( A1 => n13580, A2 => n13581, ZN => n13584);
   U6927 : INV_X1 port map( A => n13580, ZN => n13583);
   U6928 : INV_X1 port map( A => n13581, ZN => n13582);
   U6929 : AOI22_X1 port map( A1 => n10921, A2 => n13584, B1 => n13583, B2 => 
                           n13582, ZN => n13590);
   U6930 : NAND2_X1 port map( A1 => n13585, A2 => n13586, ZN => n13588);
   U6931 : XNOR2_X1 port map( A => n13588, B => n13587, ZN => n13591);
   U6932 : NAND2_X1 port map( A1 => n13590, A2 => n13591, ZN => n13596);
   U6933 : INV_X1 port map( A => n14824, ZN => n13589);
   U6934 : NAND2_X1 port map( A1 => n13596, A2 => n13589, ZN => n13594);
   U6935 : INV_X1 port map( A => n13590, ZN => n13593);
   U6936 : INV_X1 port map( A => n13591, ZN => n13592);
   U6937 : NAND2_X1 port map( A1 => n13593, A2 => n13592, ZN => n13595);
   U6938 : NAND2_X1 port map( A1 => n13594, A2 => n13595, ZN => n14863);
   U6939 : NAND2_X1 port map( A1 => n13596, A2 => n13595, ZN => n14820);
   U6940 : XNOR2_X1 port map( A => n13598, B => n13597, ZN => n13600);
   U6941 : XNOR2_X1 port map( A => n13600, B => n14965, ZN => n14862);
   U6942 : AND4_X1 port map( A1 => n10767, A2 => n10755, A3 => n10766, A4 => 
                           n10756, ZN => n14743);
   U6943 : OAI22_X1 port map( A1 => n10756, A2 => n10757, B1 => n10766, B2 => 
                           n10767, ZN => n14749);
   U6944 : INV_X1 port map( A => n14850, ZN => n14835);
   U6945 : XNOR2_X1 port map( A => n13605, B => n13604, ZN => n13615);
   U6946 : INV_X1 port map( A => n13606, ZN => n13611);
   U6947 : NAND3_X1 port map( A1 => n13609, A2 => n13608, A3 => n12410, ZN => 
                           n13610);
   U6948 : AOI21_X1 port map( B1 => n13612, B2 => n13611, A => n13610, ZN => 
                           n13614);
   U6949 : NAND2_X1 port map( A1 => n13614, A2 => n13615, ZN => n13613);
   U6950 : OAI21_X1 port map( B1 => n13615, B2 => n13614, A => n13613, ZN => 
                           n8409);
   U6951 : INV_X1 port map( A => intadd_58_n1, ZN => n13620);
   U6952 : INV_X1 port map( A => n13617, ZN => n13619);
   U6953 : NOR2_X1 port map( A1 => FP_A(0), A2 => n12567, ZN => n14585);
   U6954 : NAND2_X1 port map( A1 => n13622, A2 => n13621, ZN => n13625);
   U6955 : INV_X1 port map( A => n13623, ZN => n13624);
   U6956 : XNOR2_X1 port map( A => n13625, B => n13624, ZN => n13627);
   U6957 : XNOR2_X1 port map( A => n10828, B => n10827, ZN => n14768);
   U6958 : INV_X1 port map( A => FP_A(6), ZN => n13628);
   U6959 : XNOR2_X1 port map( A => n13628, B => n14596, ZN => n14662);
   U6960 : NAND2_X1 port map( A1 => n13630, A2 => n13629, ZN => n13633);
   U6961 : AOI22_X1 port map( A1 => n10703, A2 => n13633, B1 => n13632, B2 => 
                           n13631, ZN => n13635);
   U6962 : XNOR2_X1 port map( A => n13635, B => n13634, ZN => n13636);
   U6963 : INV_X1 port map( A => n14258, ZN => n13660);
   U6964 : INV_X1 port map( A => n13640, ZN => n13638);
   U6965 : OAI21_X1 port map( B1 => n13638, B2 => n13639, A => n13637, ZN => 
                           n13642);
   U6966 : NAND2_X1 port map( A1 => n13639, A2 => n13638, ZN => n13641);
   U6967 : NOR2_X1 port map( A1 => n13644, A2 => n13643, ZN => n13649);
   U6968 : NAND2_X1 port map( A1 => n13644, A2 => n13643, ZN => n13646);
   U6969 : NAND2_X1 port map( A1 => n13646, A2 => n13650, ZN => n13645);
   U6970 : OAI21_X1 port map( B1 => n13649, B2 => n13650, A => n13645, ZN => 
                           n13655);
   U6971 : INV_X1 port map( A => n13651, ZN => n13648);
   U6972 : NAND3_X1 port map( A1 => n13648, A2 => n13647, A3 => n13646, ZN => 
                           n13654);
   U6973 : INV_X1 port map( A => n13649, ZN => n13652);
   U6974 : NAND3_X1 port map( A1 => n13652, A2 => n13651, A3 => n13650, ZN => 
                           n13653);
   U6975 : NAND3_X1 port map( A1 => n13655, A2 => n13654, A3 => n13653, ZN => 
                           n13657);
   U6976 : XNOR2_X1 port map( A => n13657, B => n13656, ZN => n14256);
   U6977 : INV_X1 port map( A => n13663, ZN => n13664);
   U6978 : NAND2_X1 port map( A1 => n13665, A2 => n13664, ZN => n13667);
   U6979 : NAND2_X1 port map( A1 => n13667, A2 => n13666, ZN => n13672);
   U6980 : NOR2_X1 port map( A1 => n13672, A2 => n13671, ZN => n14212);
   U6981 : AND2_X1 port map( A1 => n13672, A2 => n13671, ZN => n14211);
   U6982 : NOR2_X1 port map( A1 => n14212, A2 => n14211, ZN => n13673);
   U6983 : XNOR2_X1 port map( A => n14214, B => n13673, ZN => n14869);
   U6984 : XNOR2_X1 port map( A => n13675, B => n13674, ZN => n13680);
   U6985 : XNOR2_X1 port map( A => n13677, B => n13676, ZN => n13679);
   U6986 : MUX2_X1 port map( A => n13680, B => n13679, S => n13678, Z => n14867
                           );
   U6987 : INV_X1 port map( A => n14867, ZN => n14847);
   U6988 : INV_X1 port map( A => FP_A(20), ZN => n13681);
   U6989 : XNOR2_X1 port map( A => FP_A(19), B => n13681, ZN => n14703);
   U6990 : INV_X1 port map( A => n13682, ZN => n13684);
   U6991 : INV_X1 port map( A => n13690, ZN => n13683);
   U6992 : NOR3_X1 port map( A1 => n13685, A2 => n13684, A3 => n13683, ZN => 
                           n13687);
   U6993 : AND3_X1 port map( A1 => n13688, A2 => n13687, A3 => n13686, ZN => 
                           n13699);
   U6994 : NAND2_X1 port map( A1 => n13747, A2 => n13699, ZN => n13717);
   U6995 : AOI21_X1 port map( B1 => n13691, B2 => n13690, A => n13689, ZN => 
                           n13707);
   U6996 : NAND2_X1 port map( A1 => n13717, A2 => n13707, ZN => n13692);
   U6997 : NAND3_X1 port map( A1 => n13692, A2 => n10824, A3 => n10821, ZN => 
                           n13706);
   U6998 : INV_X1 port map( A => n13699, ZN => n13697);
   U6999 : INV_X1 port map( A => n13707, ZN => n13713);
   U7000 : INV_X1 port map( A => n13709, ZN => n13693);
   U7001 : NOR2_X1 port map( A1 => n13693, A2 => n14366, ZN => n13694);
   U7002 : NOR2_X1 port map( A1 => n13713, A2 => n13694, ZN => n13700);
   U7003 : NOR2_X1 port map( A1 => n10824, A2 => n10821, ZN => n13698);
   U7004 : INV_X1 port map( A => n13698, ZN => n13695);
   U7005 : NOR2_X1 port map( A1 => n13707, A2 => n13695, ZN => n13696);
   U7006 : AOI21_X1 port map( B1 => n13697, B2 => n13700, A => n13696, ZN => 
                           n13705);
   U7007 : NAND3_X1 port map( A1 => n13747, A2 => n13699, A3 => n13698, ZN => 
                           n13704);
   U7008 : NAND3_X1 port map( A1 => n13702, A2 => n13701, A3 => n13700, ZN => 
                           n13703);
   U7009 : NAND4_X1 port map( A1 => n13706, A2 => n13705, A3 => n13704, A4 => 
                           n13703, ZN => I2_dtemp_43_port);
   U7010 : NOR2_X1 port map( A1 => n14366, A2 => n13708, ZN => n13712);
   U7011 : INV_X1 port map( A => n13712, ZN => n13716);
   U7012 : NAND4_X1 port map( A1 => n13717, A2 => n13707, A3 => n13709, A4 => 
                           n13708, ZN => n13715);
   U7013 : NAND2_X1 port map( A1 => n13708, A2 => n10821, ZN => n13710);
   U7014 : OAI22_X1 port map( A1 => n10824, A2 => n13710, B1 => n13709, B2 => 
                           n13708, ZN => n13711);
   U7015 : AOI21_X1 port map( B1 => n13713, B2 => n13712, A => n13711, ZN => 
                           n13714);
   U7016 : OAI211_X1 port map( C1 => n13717, C2 => n13716, A => n13715, B => 
                           n13714, ZN => I2_dtemp_44_port);
   U7017 : INV_X1 port map( A => n13721, ZN => n13718);
   U7018 : NOR2_X1 port map( A1 => n13718, A2 => n13719, ZN => n13722);
   U7019 : INV_X1 port map( A => n13719, ZN => n13720);
   U7020 : NAND2_X1 port map( A1 => n13725, A2 => n13724, ZN => n13726);
   U7021 : XNOR2_X1 port map( A => n13727, B => n13726, ZN => n14219);
   U7022 : XNOR2_X1 port map( A => n13728, B => n14219, ZN => n14834);
   U7023 : INV_X1 port map( A => n13728, ZN => n14837);
   U7024 : NOR2_X1 port map( A1 => FP_A(12), A2 => n14580, ZN => n14579);
   U7025 : XNOR2_X1 port map( A => n13730, B => n13729, ZN => n13735);
   U7026 : INV_X1 port map( A => n13735, ZN => n13733);
   U7027 : AND2_X1 port map( A1 => n13733, A2 => n13732, ZN => n13737);
   U7028 : INV_X1 port map( A => n13737, ZN => n13741);
   U7029 : NAND4_X1 port map( A1 => n13747, A2 => n10700, A3 => n13734, A4 => 
                           n13735, ZN => n13740);
   U7030 : INV_X1 port map( A => n10700, ZN => n13738);
   U7031 : OAI22_X1 port map( A1 => n13735, A2 => n13734, B1 => n13733, B2 => 
                           n13732, ZN => n13736);
   U7032 : AOI21_X1 port map( B1 => n13738, B2 => n13737, A => n13736, ZN => 
                           n13739);
   U7033 : OAI211_X1 port map( C1 => n13741, C2 => n13747, A => n13740, B => 
                           n13739, ZN => I2_dtemp_41_port);
   U7034 : XNOR2_X1 port map( A => n13743, B => n13742, ZN => n13748);
   U7035 : NAND3_X1 port map( A1 => n13747, A2 => n10700, A3 => n13748, ZN => 
                           n13746);
   U7036 : OR2_X1 port map( A1 => n10700, A2 => n13748, ZN => n13745);
   U7037 : OAI211_X1 port map( C1 => n13748, C2 => n13747, A => n13746, B => 
                           n13745, ZN => n14938);
   U7038 : NAND2_X1 port map( A1 => n13752, A2 => n14691, ZN => n13755);
   U7039 : NAND3_X1 port map( A1 => n14373, A2 => n13749, A3 => n14700, ZN => 
                           n13754);
   U7040 : NOR2_X1 port map( A1 => n13749, A2 => n10759, ZN => n13751);
   U7041 : OAI22_X1 port map( A1 => n13752, A2 => n14693, B1 => n10759, B2 => 
                           n14692, ZN => n13750);
   U7042 : AOI21_X1 port map( B1 => n13752, B2 => n13751, A => n13750, ZN => 
                           n13753);
   U7043 : OAI211_X1 port map( C1 => n14373, C2 => n13755, A => n13754, B => 
                           n13753, ZN => n14916);
   U7044 : NOR2_X1 port map( A1 => n13756, A2 => n13761, ZN => n13796);
   U7045 : INV_X1 port map( A => n13777, ZN => n13766);
   U7046 : INV_X1 port map( A => n13792, ZN => n13784);
   U7047 : INV_X1 port map( A => n13757, ZN => n13759);
   U7048 : NAND2_X1 port map( A1 => n13759, A2 => n13758, ZN => n13760);
   U7049 : OAI211_X1 port map( C1 => n13766, C2 => n13761, A => n13784, B => 
                           n13760, ZN => n13795);
   U7050 : INV_X1 port map( A => n13762, ZN => n13763);
   U7051 : NOR2_X1 port map( A1 => n13764, A2 => n13763, ZN => n13793);
   U7052 : INV_X1 port map( A => n13774, ZN => n13771);
   U7053 : AND4_X1 port map( A1 => n13768, A2 => n13767, A3 => n13766, A4 => 
                           n13765, ZN => n13770);
   U7054 : NAND4_X1 port map( A1 => n13772, A2 => n13771, A3 => n13770, A4 => 
                           n13769, ZN => n13783);
   U7055 : INV_X1 port map( A => n13773, ZN => n13781);
   U7056 : NOR2_X1 port map( A1 => n13774, A2 => n13777, ZN => n13780);
   U7057 : INV_X1 port map( A => n13775, ZN => n13778);
   U7058 : OAI21_X1 port map( B1 => n13778, B2 => n13777, A => n13776, ZN => 
                           n13779);
   U7059 : AOI21_X1 port map( B1 => n13781, B2 => n13780, A => n13779, ZN => 
                           n13782);
   U7060 : NAND2_X1 port map( A1 => n13783, A2 => n13782, ZN => n14335);
   U7061 : NAND2_X1 port map( A1 => n14335, A2 => n13784, ZN => n13791);
   U7062 : INV_X1 port map( A => n13785, ZN => n13789);
   U7063 : NAND2_X1 port map( A1 => n13789, A2 => n13786, ZN => n13787);
   U7064 : OAI21_X1 port map( B1 => n13789, B2 => n13788, A => n13787, ZN => 
                           n13790);
   U7065 : OAI211_X1 port map( C1 => n13793, C2 => n13792, A => n13791, B => 
                           n13790, ZN => n13794);
   U7066 : OAI21_X1 port map( B1 => n13796, B2 => n13795, A => n13794, ZN => 
                           n14934);
   U7067 : XNOR2_X1 port map( A => n13797, B => n14481, ZN => n13798);
   U7068 : XNOR2_X1 port map( A => n13799, B => n13798, ZN => n13805);
   U7069 : XOR2_X1 port map( A => n13801, B => n13800, Z => n13802);
   U7070 : XNOR2_X1 port map( A => n13803, B => n13802, ZN => n13804);
   U7071 : NOR2_X1 port map( A1 => n13805, A2 => n13804, ZN => n14292);
   U7072 : INV_X1 port map( A => n14292, ZN => n13806);
   U7073 : NAND2_X1 port map( A1 => n13805, A2 => n13804, ZN => n14290);
   U7074 : NAND2_X1 port map( A1 => n13806, A2 => n14290, ZN => n13832);
   U7075 : MUX2_X1 port map( A => n10645, B => n14840, S => n10841, Z => n13808
                           );
   U7076 : MUX2_X1 port map( A => n13442, B => n10736, S => n14459, Z => n13807
                           );
   U7077 : OAI21_X1 port map( B1 => n14121, B2 => n13808, A => n13807, ZN => 
                           n14105);
   U7078 : INV_X1 port map( A => intadd_62_A_0_port, ZN => n13812);
   U7079 : NAND2_X1 port map( A1 => n13810, A2 => n10702, ZN => n13811);
   U7080 : NAND2_X1 port map( A1 => n13812, A2 => n13811, ZN => n14103);
   U7081 : NAND2_X1 port map( A1 => n14105, A2 => n14103, ZN => n14108);
   U7082 : AND2_X1 port map( A1 => n13813, A2 => intadd_62_A_0_port, ZN => 
                           n14107);
   U7083 : INV_X1 port map( A => n14107, ZN => n13814);
   U7084 : AND2_X1 port map( A1 => n14108, A2 => n13814, ZN => n13830);
   U7085 : MUX2_X1 port map( A => n14880, B => n10886, S => n13823, Z => n13816
                           );
   U7086 : MUX2_X1 port map( A => n13819, B => n14882, S => n10631, Z => n13815
                           );
   U7087 : AND2_X1 port map( A1 => n13816, A2 => n13815, ZN => n13829);
   U7088 : MUX2_X1 port map( A => n13817, B => n10885, S => n10631, Z => n13821
                           );
   U7089 : MUX2_X1 port map( A => n13819, B => n14882, S => n8329, Z => n13820)
                           ;
   U7090 : AND2_X1 port map( A1 => n13821, A2 => n13820, ZN => n13827);
   U7091 : OR2_X1 port map( A1 => n12146, A2 => n14114, ZN => n14113);
   U7092 : NOR2_X1 port map( A1 => n13827, A2 => n14113, ZN => n13837);
   U7093 : MUX2_X1 port map( A => n12163, B => n13824, S => n13823, Z => n13825
                           );
   U7094 : AND2_X1 port map( A1 => n13826, A2 => n13825, ZN => n13840);
   U7095 : INV_X1 port map( A => n13840, ZN => n13828);
   U7096 : NAND2_X1 port map( A1 => n13827, A2 => n14113, ZN => n13838);
   U7097 : OAI21_X1 port map( B1 => n13837, B2 => n13828, A => n13838, ZN => 
                           n13835);
   U7098 : NAND2_X1 port map( A1 => n13830, A2 => n13829, ZN => n13833);
   U7099 : INV_X1 port map( A => n13833, ZN => n13831);
   U7100 : NAND2_X1 port map( A1 => n13834, A2 => n13833, ZN => n13836);
   U7101 : XNOR2_X1 port map( A => n13836, B => n13835, ZN => 
                           intadd_62_A_2_port);
   U7102 : INV_X1 port map( A => n13837, ZN => n13839);
   U7103 : NAND2_X1 port map( A1 => n13839, A2 => n13838, ZN => n13841);
   U7104 : XNOR2_X1 port map( A => n13841, B => n13840, ZN => 
                           intadd_62_B_1_port);
   U7105 : INV_X1 port map( A => n14423, ZN => n13842);
   U7106 : NAND3_X1 port map( A1 => n13844, A2 => n13843, A3 => n13842, ZN => 
                           n13846);
   U7107 : OR2_X1 port map( A1 => n14421, A2 => I1_I1_N13, ZN => n13845);
   U7108 : AOI21_X1 port map( B1 => n13846, B2 => n13845, A => n14419, ZN => 
                           I1_isZ_tab_int);
   U7109 : NAND3_X1 port map( A1 => n14663, A2 => I1_I0_N13, A3 => n14523, ZN 
                           => n14536);
   U7110 : NAND3_X1 port map( A1 => FP_A(19), A2 => n14673, A3 => FP_A(20), ZN 
                           => n14600);
   U7111 : INV_X1 port map( A => n13848, ZN => n13850);
   U7112 : NAND2_X1 port map( A1 => n13852, A2 => n13847, ZN => n13849);
   U7113 : NAND2_X1 port map( A1 => n13850, A2 => n13849, ZN => n13851);
   U7114 : OAI21_X1 port map( B1 => n13847, B2 => n13852, A => n13851, ZN => 
                           intadd_46_A_1_port);
   U7115 : MUX2_X1 port map( A => n12146, B => n11225, S => n14785, Z => n13855
                           );
   U7116 : XNOR2_X1 port map( A => n13914, B => n11226, ZN => n13853);
   U7117 : NOR2_X1 port map( A1 => n13853, A2 => n14740, ZN => n13854);
   U7118 : NOR2_X1 port map( A1 => n13855, A2 => n13854, ZN => 
                           intadd_46_B_0_port);
   U7119 : INV_X1 port map( A => n13856, ZN => n13860);
   U7120 : NAND2_X1 port map( A1 => n13858, A2 => n13857, ZN => n13859);
   U7121 : XNOR2_X1 port map( A => n13860, B => n13859, ZN => 
                           intadd_58_B_2_port);
   U7122 : XNOR2_X1 port map( A => n13862, B => n13861, ZN => n13863);
   U7123 : XNOR2_X1 port map( A => n13864, B => n13863, ZN => 
                           intadd_58_B_1_port);
   U7124 : MUX2_X1 port map( A => n13323, B => n11743, S => n14594, Z => n13865
                           );
   U7125 : INV_X1 port map( A => n13865, ZN => n13867);
   U7126 : MUX2_X1 port map( A => n10640, B => n13868, S => n10864, Z => n13866
                           );
   U7127 : NAND2_X1 port map( A1 => n13867, A2 => n13866, ZN => 
                           intadd_58_A_0_port);
   U7128 : NAND2_X1 port map( A1 => n11743, A2 => n10864, ZN => n13869);
   U7129 : NAND2_X1 port map( A1 => n13869, A2 => n13868, ZN => 
                           intadd_58_B_0_port);
   U7130 : MUX2_X1 port map( A => n14017, B => n13984, S => n10904, Z => n13871
                           );
   U7131 : MUX2_X1 port map( A => n13915, B => n14779, S => n13924, Z => n13870
                           );
   U7132 : NAND2_X1 port map( A1 => n13871, A2 => n13870, ZN => intadd_58_CI);
   U7133 : XNOR2_X1 port map( A => n13873, B => n13872, ZN => n13876);
   U7134 : INV_X1 port map( A => n13874, ZN => n13875);
   U7135 : XNOR2_X1 port map( A => n13876, B => n13875, ZN => 
                           intadd_66_A_0_port);
   U7136 : XNOR2_X1 port map( A => n13879, B => n13878, ZN => n13880);
   U7137 : XNOR2_X1 port map( A => n13877, B => n13880, ZN => 
                           intadd_66_B_0_port);
   U7138 : XNOR2_X1 port map( A => n13882, B => n13881, ZN => n13883);
   U7139 : NOR2_X1 port map( A1 => n13884, A2 => n13885, ZN => n13886);
   U7140 : NOR2_X1 port map( A1 => n11555, A2 => n13886, ZN => n13890);
   U7141 : XNOR2_X1 port map( A => n13888, B => n13887, ZN => n13889);
   U7142 : XNOR2_X1 port map( A => n13890, B => n13889, ZN => 
                           intadd_66_A_1_port);
   U7143 : XOR2_X1 port map( A => FP_B(12), B => FP_A(7), Z => n14572);
   U7144 : INV_X1 port map( A => n13891, ZN => n13892);
   U7145 : XNOR2_X1 port map( A => n13893, B => n13892, ZN => n13894);
   U7146 : FA_X1 port map( A => n13896, B => n13895, CI => n13894, CO => n14757
                           , S => n_1345);
   U7147 : OR2_X1 port map( A1 => intadd_66_SUM_1_port, A2 => n13898, ZN => 
                           n14742);
   U7148 : NAND2_X1 port map( A1 => n14742, A2 => n13897, ZN => n13900);
   U7149 : NAND2_X1 port map( A1 => n10678, A2 => n13898, ZN => n13899);
   U7150 : NAND2_X1 port map( A1 => n13900, A2 => n13899, ZN => n14754);
   U7151 : INV_X1 port map( A => n13901, ZN => n13902);
   U7152 : XNOR2_X1 port map( A => intadd_58_SUM_0_port, B => n13902, ZN => 
                           n13907);
   U7153 : INV_X1 port map( A => n13903, ZN => n13905);
   U7154 : XNOR2_X1 port map( A => n13905, B => n13904, ZN => n13906);
   U7155 : XNOR2_X1 port map( A => n13907, B => n13906, ZN => n14057);
   U7156 : MUX2_X1 port map( A => n13979, B => n13908, S => n14785, Z => n13911
                           );
   U7157 : MUX2_X1 port map( A => n13920, B => n14728, S => n14025, Z => n13909
                           );
   U7158 : INV_X1 port map( A => n13909, ZN => n13910);
   U7159 : OR2_X1 port map( A1 => n13911, A2 => n13910, ZN => n13944);
   U7160 : MUX2_X1 port map( A => n14020, B => n10939, S => n10905, Z => n13913
                           );
   U7161 : NAND2_X1 port map( A1 => n12230, A2 => n14788, ZN => n13912);
   U7162 : AND2_X1 port map( A1 => n13913, A2 => n13912, ZN => n13941);
   U7163 : XNOR2_X1 port map( A => n13944, B => n13941, ZN => n13960);
   U7164 : MUX2_X1 port map( A => n14017, B => n13984, S => n14731, Z => n13917
                           );
   U7165 : MUX2_X1 port map( A => n13915, B => n14779, S => n13914, Z => n13916
                           );
   U7166 : NAND2_X1 port map( A1 => n13917, A2 => n13916, ZN => n13958);
   U7167 : XNOR2_X1 port map( A => n13960, B => n13958, ZN => n13931);
   U7168 : OAI21_X1 port map( B1 => n13919, B2 => n13918, A => n13947, ZN => 
                           n13961);
   U7169 : NAND2_X1 port map( A1 => n13931, A2 => n13961, ZN => n13934);
   U7170 : MUX2_X1 port map( A => n13979, B => n13908, S => n14447, Z => n13928
                           );
   U7171 : MUX2_X1 port map( A => n13920, B => n14728, S => n14594, Z => n13923
                           );
   U7172 : INV_X1 port map( A => n13923, ZN => n13921);
   U7173 : OR2_X1 port map( A1 => n13928, A2 => n13921, ZN => n13988);
   U7174 : NAND2_X1 port map( A1 => n13988, A2 => n13922, ZN => n13930);
   U7175 : NAND2_X1 port map( A1 => n13923, A2 => n13965, ZN => n13927);
   U7176 : MUX2_X1 port map( A => n14020, B => n10940, S => n13924, Z => n13926
                           );
   U7177 : NAND2_X1 port map( A1 => n12230, A2 => n14448, ZN => n13925);
   U7178 : NAND2_X1 port map( A1 => n13926, A2 => n13925, ZN => n13966);
   U7179 : OAI21_X1 port map( B1 => n13928, B2 => n13927, A => n13966, ZN => 
                           n13929);
   U7180 : NAND2_X1 port map( A1 => n13930, A2 => n13929, ZN => n13959);
   U7181 : INV_X1 port map( A => n13931, ZN => n13933);
   U7182 : INV_X1 port map( A => n13961, ZN => n13932);
   U7183 : AOI22_X1 port map( A1 => n13934, A2 => n13959, B1 => n13933, B2 => 
                           n13932, ZN => n13978);
   U7184 : XNOR2_X1 port map( A => n13936, B => n13935, ZN => n13948);
   U7185 : XNOR2_X1 port map( A => n13938, B => n13937, ZN => n13939);
   U7186 : XNOR2_X1 port map( A => n13940, B => n13939, ZN => n13950);
   U7187 : XNOR2_X1 port map( A => n13948, B => n13950, ZN => n13946);
   U7188 : INV_X1 port map( A => n13941, ZN => n13942);
   U7189 : AND2_X1 port map( A1 => n13958, A2 => n13942, ZN => n13943);
   U7190 : OAI22_X1 port map( A1 => n13944, A2 => n13943, B1 => n13958, B2 => 
                           n13942, ZN => n13949);
   U7191 : XNOR2_X1 port map( A => n13949, B => n13947, ZN => n13945);
   U7192 : XNOR2_X1 port map( A => n13946, B => n13945, ZN => n13977);
   U7193 : XNOR2_X1 port map( A => n13948, B => n13947, ZN => n13951);
   U7194 : OAI21_X1 port map( B1 => n13951, B2 => n13950, A => n13949, ZN => 
                           n13953);
   U7195 : NAND2_X1 port map( A1 => n13951, A2 => n13950, ZN => n13952);
   U7196 : NAND2_X1 port map( A1 => n13953, A2 => n13952, ZN => n13957);
   U7197 : OAI21_X1 port map( B1 => n13978, B2 => n13977, A => n13957, ZN => 
                           n13956);
   U7198 : NOR2_X1 port map( A1 => n13978, A2 => n13957, ZN => n13955);
   U7199 : INV_X1 port map( A => n13977, ZN => n13954);
   U7200 : AOI22_X1 port map( A1 => n14057, A2 => n13956, B1 => n13955, B2 => 
                           n13954, ZN => n14061);
   U7201 : INV_X1 port map( A => n13957, ZN => n14056);
   U7202 : XNOR2_X1 port map( A => n13959, B => n13958, ZN => n13964);
   U7203 : INV_X1 port map( A => n13960, ZN => n13962);
   U7204 : XNOR2_X1 port map( A => n13962, B => n13961, ZN => n13963);
   U7205 : XNOR2_X1 port map( A => n13964, B => n13963, ZN => n14053);
   U7206 : XNOR2_X1 port map( A => n13966, B => n13965, ZN => n13989);
   U7207 : XNOR2_X1 port map( A => n13988, B => n13989, ZN => n13973);
   U7208 : AOI21_X1 port map( B1 => n10938, B2 => n14719, A => n13968, ZN => 
                           n13995);
   U7209 : MUX2_X1 port map( A => n14020, B => n10940, S => n8401, Z => n13970)
                           ;
   U7210 : NAND2_X1 port map( A1 => n14771, A2 => n14465, ZN => n13969);
   U7211 : NAND2_X1 port map( A1 => n13970, A2 => n13969, ZN => n13994);
   U7212 : NAND2_X1 port map( A1 => n13995, A2 => n13994, ZN => n13974);
   U7213 : NAND2_X1 port map( A1 => n13973, A2 => n13974, ZN => n13976);
   U7214 : MUX2_X1 port map( A => n14017, B => n13984, S => n13914, Z => n13972
                           );
   U7215 : MUX2_X1 port map( A => n14779, B => n14456, S => n14593, Z => n13971
                           );
   U7216 : NAND2_X1 port map( A1 => n13972, A2 => n13971, ZN => n13990);
   U7217 : INV_X1 port map( A => n13973, ZN => n13975);
   U7218 : INV_X1 port map( A => n13974, ZN => n13987);
   U7219 : AOI22_X1 port map( A1 => n13976, A2 => n13990, B1 => n13975, B2 => 
                           n13987, ZN => n14052);
   U7220 : AOI22_X1 port map( A1 => n13978, A2 => n13977, B1 => n14053, B2 => 
                           n14052, ZN => n14055);
   U7221 : MUX2_X1 port map( A => n13979, B => n13908, S => n14777, Z => n13983
                           );
   U7222 : MUX2_X1 port map( A => n13920, B => n14728, S => n10864, Z => n13981
                           );
   U7223 : INV_X1 port map( A => n13981, ZN => n13982);
   U7224 : OR2_X1 port map( A1 => n13983, A2 => n13982, ZN => n14011);
   U7225 : MUX2_X1 port map( A => n11201, B => n14017, S => n14593, Z => n13986
                           );
   U7226 : MUX2_X1 port map( A => n14779, B => n14456, S => n14025, Z => n13985
                           );
   U7227 : AND2_X1 port map( A1 => n13986, A2 => n13985, ZN => n13997);
   U7228 : INV_X1 port map( A => n13997, ZN => n14010);
   U7229 : NAND2_X1 port map( A1 => n14011, A2 => n14010, ZN => n14012);
   U7230 : INV_X1 port map( A => n14012, ZN => n14007);
   U7231 : XNOR2_X1 port map( A => n13988, B => n13987, ZN => n13993);
   U7232 : INV_X1 port map( A => n13989, ZN => n13991);
   U7233 : XNOR2_X1 port map( A => n13991, B => n13990, ZN => n13992);
   U7234 : XNOR2_X1 port map( A => n13995, B => n13994, ZN => n14008);
   U7235 : NAND2_X1 port map( A1 => n13997, A2 => n14008, ZN => n13996);
   U7236 : XNOR2_X1 port map( A => n14011, B => n13996, ZN => n13999);
   U7237 : NOR2_X1 port map( A1 => n14008, A2 => n13997, ZN => n13998);
   U7238 : OAI22_X1 port map( A1 => n13999, A2 => n13998, B1 => n14012, B2 => 
                           n14008, ZN => n14049);
   U7239 : MUX2_X1 port map( A => n13984, B => n14017, S => n14025, Z => n14001
                           );
   U7240 : MUX2_X1 port map( A => n14779, B => n14456, S => n14594, Z => n14000
                           );
   U7241 : NAND2_X1 port map( A1 => n14001, A2 => n14000, ZN => n14031);
   U7242 : AND2_X1 port map( A1 => n14002, A2 => n14719, ZN => n14028);
   U7243 : MUX2_X1 port map( A => n14020, B => n10939, S => n10635, Z => n14004
                           );
   U7244 : NAND2_X1 port map( A1 => n12230, A2 => n14593, ZN => n14003);
   U7245 : NAND2_X1 port map( A1 => n14004, A2 => n14003, ZN => n14029);
   U7246 : OAI21_X1 port map( B1 => n14031, B2 => n14028, A => n14029, ZN => 
                           n14006);
   U7247 : NAND2_X1 port map( A1 => n14031, A2 => n14028, ZN => n14005);
   U7248 : NAND2_X1 port map( A1 => n14006, A2 => n14005, ZN => n14048);
   U7249 : OAI211_X1 port map( C1 => n14007, C2 => n14045, A => n14049, B => 
                           n14048, ZN => n14015);
   U7250 : INV_X1 port map( A => n14008, ZN => n14009);
   U7251 : OAI21_X1 port map( B1 => n14011, B2 => n14010, A => n14009, ZN => 
                           n14013);
   U7252 : NAND2_X1 port map( A1 => n14013, A2 => n14012, ZN => n14046);
   U7253 : NAND2_X1 port map( A1 => n14045, A2 => n14046, ZN => n14014);
   U7254 : AND2_X1 port map( A1 => n14015, A2 => n14014, ZN => n14051);
   U7255 : INV_X1 port map( A => n14017, ZN => n14016);
   U7256 : AOI21_X1 port map( B1 => n14016, B2 => n10864, A => n14484, ZN => 
                           n14033);
   U7257 : MUX2_X1 port map( A => n11201, B => n14017, S => n14594, Z => n14035
                           );
   U7258 : MUX2_X1 port map( A => n10940, B => n14020, S => n14593, Z => n14019
                           );
   U7259 : NAND2_X1 port map( A1 => n14771, A2 => n14025, ZN => n14018);
   U7260 : AND2_X1 port map( A1 => n14019, A2 => n14018, ZN => n14036);
   U7261 : NAND2_X1 port map( A1 => n12230, A2 => n14594, ZN => n14023);
   U7262 : MUX2_X1 port map( A => n10940, B => n14020, S => n14025, Z => n14022
                           );
   U7263 : AOI21_X1 port map( B1 => n14023, B2 => n14022, A => n14499, ZN => 
                           n14024);
   U7264 : OAI21_X1 port map( B1 => n14035, B2 => n14036, A => n14024, ZN => 
                           n14027);
   U7265 : NAND3_X1 port map( A1 => n14784, A2 => n14594, A3 => n14025, ZN => 
                           n14026);
   U7266 : MUX2_X1 port map( A => n14027, B => n14026, S => n10864, Z => n14039
                           );
   U7267 : INV_X1 port map( A => n14028, ZN => n14030);
   U7268 : XNOR2_X1 port map( A => n14030, B => n14029, ZN => n14032);
   U7269 : XNOR2_X1 port map( A => n14032, B => n14031, ZN => n14038);
   U7270 : AOI21_X1 port map( B1 => n14033, B2 => n14039, A => n14038, ZN => 
                           n14043);
   U7271 : MUX2_X1 port map( A => n14779, B => n14456, S => n10864, Z => n14034
                           );
   U7272 : NAND2_X1 port map( A1 => n14035, A2 => n14034, ZN => n14040);
   U7273 : INV_X1 port map( A => n14036, ZN => n14041);
   U7274 : NAND2_X1 port map( A1 => n14040, A2 => n14041, ZN => n14037);
   U7275 : AOI21_X1 port map( B1 => n14039, B2 => n14038, A => n14037, ZN => 
                           n14042);
   U7276 : OAI22_X1 port map( A1 => n14043, A2 => n14042, B1 => n14041, B2 => 
                           n14040, ZN => n14044);
   U7277 : INV_X1 port map( A => n14044, ZN => n14047);
   U7278 : OAI211_X1 port map( C1 => n14053, C2 => n14052, A => n14051, B => 
                           n14050, ZN => n14054);
   U7279 : OAI211_X1 port map( C1 => n14057, C2 => n14056, A => n14055, B => 
                           n14054, ZN => n14060);
   U7280 : AOI22_X1 port map( A1 => n14061, A2 => n14060, B1 => n14059, B2 => 
                           n14058, ZN => n14746);
   U7281 : XNOR2_X1 port map( A => n14062, B => intadd_46_SUM_1_port, ZN => 
                           n14064);
   U7282 : INV_X1 port map( A => n14066, ZN => n14063);
   U7283 : XNOR2_X1 port map( A => n14064, B => n14063, ZN => n14761);
   U7284 : INV_X1 port map( A => intadd_66_n1, ZN => n14767);
   U7285 : XNOR2_X1 port map( A => n14065, B => intadd_46_SUM_1_port, ZN => 
                           n14067);
   U7286 : XNOR2_X1 port map( A => n14067, B => n10687, ZN => n14773);
   U7287 : NAND2_X1 port map( A1 => n14069, A2 => n14068, ZN => n14072);
   U7288 : INV_X1 port map( A => n14070, ZN => n14071);
   U7289 : XNOR2_X1 port map( A => n14072, B => n14071, ZN => n14800);
   U7290 : NAND2_X1 port map( A1 => n14073, A2 => n14074, ZN => n14076);
   U7291 : XNOR2_X1 port map( A => n14076, B => n14075, ZN => 
                           intadd_46_B_4_port);
   U7292 : INV_X1 port map( A => n14801, ZN => n14077);
   U7293 : NOR2_X1 port map( A1 => n14077, A2 => n14800, ZN => n14797);
   U7294 : NAND2_X1 port map( A1 => n14077, A2 => n14800, ZN => n14798);
   U7295 : FA_X1 port map( A => n10918, B => n14189, CI => n14188, CO => n14082
                           , S => n_1346);
   U7296 : XNOR2_X1 port map( A => n14079, B => n14078, ZN => n14080);
   U7297 : XNOR2_X1 port map( A => n14081, B => n14080, ZN => n14194);
   U7298 : XNOR2_X1 port map( A => n14082, B => n14194, ZN => n14806);
   U7299 : OAI21_X1 port map( B1 => n14085, B2 => n14083, A => n14084, ZN => 
                           n14091);
   U7300 : INV_X1 port map( A => n14086, ZN => n14089);
   U7301 : OAI211_X1 port map( C1 => n14089, C2 => n14088, A => n14087, B => 
                           n14083, ZN => n14090);
   U7302 : NAND2_X1 port map( A1 => n14091, A2 => n14090, ZN => n14816);
   U7303 : NAND2_X1 port map( A1 => n14093, A2 => n14092, ZN => n14096);
   U7304 : NAND3_X1 port map( A1 => n14096, A2 => n14095, A3 => n14094, ZN => 
                           n14790);
   U7305 : INV_X1 port map( A => n14097, ZN => n14812);
   U7306 : NAND2_X1 port map( A1 => n14099, A2 => n14098, ZN => n14102);
   U7307 : INV_X1 port map( A => n14100, ZN => n14101);
   U7308 : NAND3_X1 port map( A1 => n10844, A2 => n10843, A3 => n10780, ZN => 
                           n14831);
   U7309 : INV_X1 port map( A => n14103, ZN => n14104);
   U7310 : NOR2_X1 port map( A1 => n14104, A2 => n14107, ZN => n14106);
   U7311 : OAI22_X1 port map( A1 => n14108, A2 => n14107, B1 => n14106, B2 => 
                           n14105, ZN => intadd_62_A_1_port);
   U7312 : XNOR2_X1 port map( A => n14110, B => n14109, ZN => n14112);
   U7313 : XNOR2_X1 port map( A => n14112, B => n14111, ZN => 
                           intadd_62_B_2_port);
   U7314 : INV_X1 port map( A => n14113, ZN => n14116);
   U7315 : NOR2_X1 port map( A1 => n14114, A2 => n11225, ZN => n14115);
   U7316 : MUX2_X1 port map( A => n14116, B => n14115, S => n14881, Z => 
                           intadd_62_B_0_port);
   U7317 : MUX2_X1 port map( A => n14840, B => n10645, S => n13261, Z => n14120
                           );
   U7318 : MUX2_X1 port map( A => n10925, B => n10736, S => n14467, Z => n14119
                           );
   U7319 : OAI21_X1 port map( B1 => n14121, B2 => n14120, A => n14119, ZN => 
                           n14122);
   U7320 : INV_X1 port map( A => n14122, ZN => intadd_62_CI);
   U7321 : INV_X1 port map( A => n14123, ZN => n14128);
   U7322 : INV_X1 port map( A => n14124, ZN => n14126);
   U7323 : NAND2_X1 port map( A1 => n14126, A2 => n14125, ZN => n14127);
   U7324 : XNOR2_X1 port map( A => n14128, B => n14127, ZN => n14278);
   U7325 : XNOR2_X1 port map( A => n14130, B => n14129, ZN => n14132);
   U7326 : INV_X1 port map( A => n14132, ZN => n14133);
   U7327 : MUX2_X1 port map( A => n14133, B => n14132, S => n14131, Z => n14276
                           );
   U7328 : XNOR2_X1 port map( A => n14278, B => n14276, ZN => n14156);
   U7329 : INV_X1 port map( A => n14134, ZN => n14136);
   U7330 : OAI21_X1 port map( B1 => n14136, B2 => n14137, A => n14135, ZN => 
                           n14139);
   U7331 : NAND2_X1 port map( A1 => n14137, A2 => n14136, ZN => n14138);
   U7332 : NAND2_X1 port map( A1 => n14139, A2 => n14138, ZN => n14267);
   U7333 : INV_X1 port map( A => n14267, ZN => n14153);
   U7334 : INV_X1 port map( A => n14143, ZN => n14141);
   U7335 : NAND2_X1 port map( A1 => n14141, A2 => n14140, ZN => n14148);
   U7336 : NAND2_X1 port map( A1 => n14143, A2 => n14142, ZN => n14146);
   U7337 : INV_X1 port map( A => n14144, ZN => n14145);
   U7338 : NAND2_X1 port map( A1 => n14146, A2 => n14145, ZN => n14147);
   U7339 : NAND2_X1 port map( A1 => n14148, A2 => n14147, ZN => n14271);
   U7340 : AND2_X1 port map( A1 => n14153, A2 => n14271, ZN => n14154);
   U7341 : XNOR2_X1 port map( A => n14150, B => n14149, ZN => n14152);
   U7342 : XNOR2_X1 port map( A => n14152, B => n14151, ZN => n14270);
   U7343 : OAI22_X1 port map( A1 => n14154, A2 => n14270, B1 => n14153, B2 => 
                           n14271, ZN => n14155);
   U7344 : XNOR2_X1 port map( A => n14156, B => n14155, ZN => 
                           intadd_42_A_3_port);
   U7345 : XNOR2_X1 port map( A => n14158, B => n14157, ZN => n14160);
   U7346 : XNOR2_X1 port map( A => n14160, B => n14159, ZN => 
                           intadd_42_B_3_port);
   U7347 : XNOR2_X1 port map( A => n14162, B => n14161, ZN => n14164);
   U7348 : XNOR2_X1 port map( A => n14164, B => n14163, ZN => n14179);
   U7349 : INV_X1 port map( A => n14179, ZN => n14175);
   U7350 : INV_X1 port map( A => n14171, ZN => n14166);
   U7351 : INV_X1 port map( A => n14170, ZN => n14165);
   U7352 : NAND2_X1 port map( A1 => n14166, A2 => n14165, ZN => n14167);
   U7353 : NAND3_X1 port map( A1 => n14169, A2 => n14168, A3 => n14167, ZN => 
                           n14173);
   U7354 : NAND2_X1 port map( A1 => n14171, A2 => n14170, ZN => n14172);
   U7355 : AND2_X1 port map( A1 => n14173, A2 => n14172, ZN => n14180);
   U7356 : INV_X1 port map( A => n14180, ZN => n14174);
   U7357 : NAND2_X1 port map( A1 => n14175, A2 => n14174, ZN => n14240);
   U7358 : INV_X1 port map( A => n14240, ZN => n14182);
   U7359 : NAND2_X1 port map( A1 => n14177, A2 => n14176, ZN => n14239);
   U7360 : INV_X1 port map( A => n14238, ZN => n14178);
   U7361 : NAND2_X1 port map( A1 => n14178, A2 => n14240, ZN => n14181);
   U7362 : NAND2_X1 port map( A1 => n14180, A2 => n14179, ZN => n14241);
   U7363 : OAI211_X1 port map( C1 => n14182, C2 => n14239, A => n14181, B => 
                           n14241, ZN => intadd_42_n11);
   U7364 : INV_X1 port map( A => n10686, ZN => n14183);
   U7365 : NAND2_X1 port map( A1 => n14183, A2 => intadd_46_SUM_2_port, ZN => 
                           n14795);
   U7366 : INV_X1 port map( A => intadd_46_SUM_2_port, ZN => n14184);
   U7367 : NAND2_X1 port map( A1 => n14184, A2 => n14796, ZN => n14799);
   U7369 : XNOR2_X1 port map( A => n14816, B => n14963, ZN => n14186);
   U7370 : XNOR2_X1 port map( A => n14186, B => n14185, ZN => n14808);
   U7371 : INV_X1 port map( A => n14187, ZN => n14814);
   U7372 : AOI21_X1 port map( B1 => n14190, B2 => n14189, A => n14188, ZN => 
                           n14192);
   U7373 : NOR2_X1 port map( A1 => n14190, A2 => n14189, ZN => n14191);
   U7374 : NOR2_X1 port map( A1 => n14192, A2 => n14191, ZN => n14195);
   U7375 : NAND2_X1 port map( A1 => n14195, A2 => n14194, ZN => n14193);
   U7376 : NAND2_X1 port map( A1 => n14193, A2 => n14816, ZN => n14198);
   U7377 : INV_X1 port map( A => n14194, ZN => n14196);
   U7378 : NAND2_X1 port map( A1 => n14196, A2 => n10917, ZN => n14197);
   U7379 : NAND2_X1 port map( A1 => n14198, A2 => n14197, ZN => n14817);
   U7380 : INV_X1 port map( A => n14197, ZN => n14821);
   U7381 : INV_X1 port map( A => n14198, ZN => n14822);
   U7382 : XNOR2_X1 port map( A => n14199, B => n14862, ZN => n14826);
   U7383 : INV_X1 port map( A => n14829, ZN => n14210);
   U7384 : INV_X1 port map( A => n14200, ZN => n14209);
   U7385 : OAI21_X1 port map( B1 => n14963, B2 => n13550, A => n14202, ZN => 
                           n14205);
   U7387 : INV_X1 port map( A => n14211, ZN => n14213);
   U7388 : AOI21_X1 port map( B1 => n14214, B2 => n14213, A => n14212, ZN => 
                           n14849);
   U7389 : NAND2_X1 port map( A1 => n14216, A2 => n14215, ZN => n14218);
   U7390 : XNOR2_X1 port map( A => n14218, B => n14217, ZN => n14848);
   U7391 : INV_X1 port map( A => n14848, ZN => n14836);
   U7392 : INV_X1 port map( A => n14219, ZN => n14838);
   U7393 : NAND2_X1 port map( A1 => n14221, A2 => n14220, ZN => n14223);
   U7394 : NAND2_X1 port map( A1 => n14223, A2 => n14222, ZN => n14249);
   U7395 : NAND2_X1 port map( A1 => n14225, A2 => n14224, ZN => n14227);
   U7396 : XNOR2_X1 port map( A => n14227, B => n14226, ZN => n14250);
   U7397 : XNOR2_X1 port map( A => n14249, B => n14250, ZN => n14843);
   U7398 : NAND2_X1 port map( A1 => n14229, A2 => n14228, ZN => n14231);
   U7399 : XNOR2_X1 port map( A => n14231, B => n14230, ZN => n14854);
   U7400 : INV_X1 port map( A => n14232, ZN => n14233);
   U7401 : NAND2_X1 port map( A1 => n14234, A2 => n14233, ZN => n14236);
   U7402 : NAND2_X1 port map( A1 => n14236, A2 => n14235, ZN => n14245);
   U7403 : XNOR2_X1 port map( A => n14271, B => n14267, ZN => n14237);
   U7404 : XNOR2_X1 port map( A => n14237, B => n14270, ZN => n14244);
   U7405 : XNOR2_X1 port map( A => n14245, B => n14244, ZN => n14851);
   U7406 : NAND2_X1 port map( A1 => n14239, A2 => n14238, ZN => n14243);
   U7407 : NAND2_X1 port map( A1 => n14241, A2 => n14240, ZN => n14242);
   U7408 : XNOR2_X1 port map( A => n14243, B => n14242, ZN => n14853);
   U7409 : OR2_X1 port map( A1 => n14252, A2 => n14251, ZN => n14872);
   U7410 : INV_X1 port map( A => n14244, ZN => n14246);
   U7411 : OAI21_X1 port map( B1 => n14853, B2 => n14246, A => n14245, ZN => 
                           n14248);
   U7412 : NAND2_X1 port map( A1 => n14853, A2 => n14246, ZN => n14247);
   U7413 : NAND2_X1 port map( A1 => n14248, A2 => n14247, ZN => n14897);
   U7414 : INV_X1 port map( A => n14249, ZN => n14856);
   U7415 : INV_X1 port map( A => n14250, ZN => n14855);
   U7416 : XNOR2_X1 port map( A => n14252, B => n14251, ZN => n14857);
   U7417 : NAND2_X1 port map( A1 => n11676, A2 => n14253, ZN => n14255);
   U7418 : NAND2_X1 port map( A1 => n14255, A2 => n14254, ZN => n14866);
   U7419 : XNOR2_X1 port map( A => n14257, B => n14256, ZN => n14259);
   U7420 : XNOR2_X1 port map( A => n14259, B => n14258, ZN => n14864);
   U7421 : INV_X1 port map( A => n14862, ZN => n14860);
   U7422 : INV_X1 port map( A => n14864, ZN => n14865);
   U7423 : NAND2_X1 port map( A1 => n14261, A2 => n14260, ZN => n14263);
   U7424 : XNOR2_X1 port map( A => n14263, B => n14262, ZN => n14876);
   U7425 : FA_X1 port map( A => n14266, B => n14265, CI => n14264, CO => 
                           intadd_61_n7, S => n14286);
   U7426 : NAND2_X1 port map( A1 => n14270, A2 => n14271, ZN => n14268);
   U7427 : NAND2_X1 port map( A1 => n14268, A2 => n14267, ZN => n14269);
   U7428 : OAI21_X1 port map( B1 => n14271, B2 => n14270, A => n14269, ZN => 
                           n14282);
   U7429 : INV_X1 port map( A => n14278, ZN => n14272);
   U7430 : OAI21_X1 port map( B1 => n14282, B2 => n14272, A => n14276, ZN => 
                           n14274);
   U7431 : NAND2_X1 port map( A1 => n14282, A2 => n14272, ZN => n14273);
   U7432 : AND2_X1 port map( A1 => n14274, A2 => n14273, ZN => n14275);
   U7433 : OR2_X1 port map( A1 => n14286, A2 => n14275, ZN => n14874);
   U7434 : NAND2_X1 port map( A1 => n14286, A2 => n14275, ZN => n14875);
   U7435 : INV_X1 port map( A => n14286, ZN => n14277);
   U7436 : INV_X1 port map( A => n14276, ZN => n14279);
   U7437 : NAND2_X1 port map( A1 => n14279, A2 => n14278, ZN => n14280);
   U7438 : NAND3_X1 port map( A1 => n14277, A2 => n14282, A3 => n14280, ZN => 
                           n14289);
   U7439 : NOR2_X1 port map( A1 => n14279, A2 => n14278, ZN => n14283);
   U7440 : NAND2_X1 port map( A1 => n14286, A2 => n14280, ZN => n14281);
   U7441 : OAI21_X1 port map( B1 => n14286, B2 => n14283, A => n14281, ZN => 
                           n14288);
   U7442 : INV_X1 port map( A => n14282, ZN => n14285);
   U7443 : INV_X1 port map( A => n14283, ZN => n14284);
   U7444 : NAND3_X1 port map( A1 => n14286, A2 => n14285, A3 => n14284, ZN => 
                           n14287);
   U7445 : NAND3_X1 port map( A1 => n14289, A2 => n14288, A3 => n14287, ZN => 
                           n14877);
   U7446 : OAI21_X1 port map( B1 => n14292, B2 => n14291, A => n14290, ZN => 
                           n14362);
   U7447 : NAND2_X1 port map( A1 => n14294, A2 => n14293, ZN => n14295);
   U7448 : XNOR2_X1 port map( A => n14296, B => n14295, ZN => n14360);
   U7449 : AND2_X1 port map( A1 => n14362, A2 => n14360, ZN => n14905);
   U7450 : NOR2_X1 port map( A1 => n14362, A2 => n14360, ZN => n14903);
   U7451 : NOR2_X1 port map( A1 => n14358, A2 => n14356, ZN => n14297);
   U7452 : NOR2_X1 port map( A1 => n14903, A2 => n14297, ZN => n14879);
   U7453 : NAND2_X1 port map( A1 => n14307, A2 => n14298, ZN => n14299);
   U7454 : MUX2_X1 port map( A => n14300, B => n14299, S => n14308, Z => n14312
                           );
   U7455 : AOI21_X1 port map( B1 => n14305, B2 => n14306, A => n14312, ZN => 
                           n14886);
   U7456 : INV_X1 port map( A => n14306, ZN => n14304);
   U7457 : INV_X1 port map( A => n14312, ZN => n14303);
   U7458 : AOI21_X1 port map( B1 => n14304, B2 => n14302, A => n14303, ZN => 
                           n14301);
   U7459 : AND2_X1 port map( A1 => n14913, A2 => n14301, ZN => n14885);
   U7460 : INV_X1 port map( A => n14885, ZN => n14884);
   U7461 : INV_X1 port map( A => n14913, ZN => n14317);
   U7462 : NAND3_X1 port map( A1 => n14304, A2 => n14303, A3 => n14302, ZN => 
                           n14315);
   U7463 : NAND3_X1 port map( A1 => n14306, A2 => n14305, A3 => n14312, ZN => 
                           n14314);
   U7464 : INV_X1 port map( A => n14307, ZN => n14311);
   U7465 : NAND2_X1 port map( A1 => n14309, A2 => n14308, ZN => n14310);
   U7466 : NAND3_X1 port map( A1 => n14312, A2 => n14311, A3 => n14310, ZN => 
                           n14313);
   U7467 : NAND3_X1 port map( A1 => n14315, A2 => n14314, A3 => n14313, ZN => 
                           n14316);
   U7468 : AOI21_X1 port map( B1 => n14317, B2 => n14886, A => n14316, ZN => 
                           n14889);
   U7469 : NAND2_X1 port map( A1 => n14319, A2 => n14318, ZN => n14320);
   U7470 : XNOR2_X1 port map( A => n14321, B => n14320, ZN => n14325);
   U7471 : MUX2_X1 port map( A => n14322, B => n14325, S => n10927, Z => n14607
                           );
   U7472 : INV_X1 port map( A => n14490, ZN => n14324);
   U7473 : MUX2_X1 port map( A => n14325, B => n14324, S => n10927, Z => n14581
                           );
   U7474 : MUX2_X1 port map( A => n14519, B => n2606, S => n10975, Z => n14327)
                           ;
   U7475 : INV_X1 port map( A => n14327, ZN => n14326);
   U7476 : XNOR2_X1 port map( A => n14328, B => n14326, ZN => I3_SIG_out_8_port
                           );
   U7477 : OR2_X1 port map( A1 => n14328, A2 => n14327, ZN => n14330);
   U7478 : MUX2_X1 port map( A => n8381, B => n8371, S => n14729, Z => n14329);
   U7479 : XNOR2_X1 port map( A => n14330, B => n14329, ZN => I3_SIG_out_9_port
                           );
   U7480 : INV_X1 port map( A => n14331, ZN => n14332);
   U7481 : XNOR2_X1 port map( A => n12248, B => n14332, ZN => 
                           I3_SIG_out_11_port);
   U7482 : XOR2_X1 port map( A => n14334, B => n14333, Z => n14337);
   U7483 : INV_X1 port map( A => n14337, ZN => n14336);
   U7484 : MUX2_X1 port map( A => n14337, B => n14336, S => n14335, Z => 
                           I2_dtemp_34_port);
   U7485 : XNOR2_X1 port map( A => n14338, B => n14340, ZN => 
                           I3_SIG_out_13_port);
   U7486 : INV_X1 port map( A => n14338, ZN => n14341);
   U7487 : AOI21_X1 port map( B1 => n14341, B2 => n14340, A => n14339, ZN => 
                           n14342);
   U7488 : NOR2_X1 port map( A1 => n14342, A2 => n14345, ZN => 
                           I3_SIG_out_14_port);
   U7489 : INV_X1 port map( A => n14343, ZN => n14344);
   U7490 : XNOR2_X1 port map( A => n14345, B => n14344, ZN => 
                           I3_SIG_out_15_port);
   U7491 : XNOR2_X1 port map( A => n14346, B => n14348, ZN => 
                           I3_SIG_out_17_port);
   U7492 : INV_X1 port map( A => n14346, ZN => n14349);
   U7493 : AOI21_X1 port map( B1 => n14349, B2 => n14348, A => n14347, ZN => 
                           n14350);
   U7494 : NOR2_X1 port map( A1 => n14350, A2 => n14353, ZN => 
                           I3_SIG_out_18_port);
   U7495 : INV_X1 port map( A => n14351, ZN => n14352);
   U7496 : XNOR2_X1 port map( A => n14353, B => n14352, ZN => 
                           I3_SIG_out_19_port);
   U7497 : NAND2_X1 port map( A1 => n14355, A2 => n14354, ZN => n14898);
   U7498 : MUX2_X1 port map( A => n14516, B => n8347, S => n14729, Z => n14901)
                           ;
   U7499 : INV_X1 port map( A => n14356, ZN => n14357);
   U7500 : XNOR2_X1 port map( A => n14358, B => n14357, ZN => n14906);
   U7501 : INV_X1 port map( A => n14903, ZN => n14904);
   U7502 : NOR2_X1 port map( A1 => n14905, A2 => n14906, ZN => n14908);
   U7503 : INV_X1 port map( A => n14362, ZN => n14363);
   U7504 : INV_X1 port map( A => n14360, ZN => n14359);
   U7505 : NAND2_X1 port map( A1 => n14906, A2 => n14360, ZN => n14361);
   U7506 : INV_X1 port map( A => n14364, ZN => n14372);
   U7507 : NAND2_X1 port map( A1 => n14373, A2 => n14372, ZN => n14369);
   U7508 : INV_X1 port map( A => n14365, ZN => n14367);
   U7509 : AOI21_X1 port map( B1 => n14368, B2 => n14367, A => n14366, ZN => 
                           n14370);
   U7510 : NAND4_X1 port map( A1 => n14369, A2 => n14370, A3 => n14707, A4 => 
                           n14706, ZN => n14376);
   U7511 : INV_X1 port map( A => n14370, ZN => n14371);
   U7512 : AOI21_X1 port map( B1 => n14371, B2 => n10788, A => n14688, ZN => 
                           n14375);
   U7513 : NAND3_X1 port map( A1 => n14373, A2 => n14372, A3 => n10788, ZN => 
                           n14374);
   U7514 : NAND3_X1 port map( A1 => n14376, A2 => n14375, A3 => n14374, ZN => 
                           n14935);
   U7515 : MUX2_X1 port map( A => n2590, B => n2589, S => SIG_in_27_port, Z => 
                           n14910);
   U7516 : INV_X1 port map( A => n14914, ZN => n14911);
   U7517 : AND2_X1 port map( A1 => n14913, A2 => n14914, ZN => n14912);
   U7518 : INV_X1 port map( A => n14912, ZN => n14915);
   U7519 : NAND2_X1 port map( A1 => n14470, A2 => n14500, ZN => n14917);
   U7520 : NAND4_X1 port map( A1 => B_EXP_2_port, A2 => B_EXP_3_port, A3 => 
                           B_EXP_4_port, A4 => B_EXP_5_port, ZN => n14379);
   U7521 : NAND3_X1 port map( A1 => B_EXP_1_port, A2 => B_EXP_6_port, A3 => 
                           B_EXP_0_port, ZN => n14378);
   U7522 : NOR2_X1 port map( A1 => B_EXP_7_port, A2 => A_EXP_7_port, ZN => 
                           n14377);
   U7523 : OAI21_X1 port map( B1 => n14379, B2 => n14378, A => n14377, ZN => 
                           n14383);
   U7524 : NAND4_X1 port map( A1 => A_EXP_2_port, A2 => A_EXP_3_port, A3 => 
                           A_EXP_4_port, A4 => A_EXP_5_port, ZN => n14381);
   U7525 : NAND3_X1 port map( A1 => A_EXP_1_port, A2 => A_EXP_6_port, A3 => 
                           A_EXP_0_port, ZN => n14380);
   U7526 : NOR2_X1 port map( A1 => n14381, A2 => n14380, ZN => n14382);
   U7527 : NOR2_X1 port map( A1 => n14383, A2 => n14382, ZN => I2_N0);
   U7528 : NOR2_X1 port map( A1 => A_EXP_1_port, A2 => B_EXP_1_port, ZN => 
                           n14385);
   U7529 : NAND2_X1 port map( A1 => B_EXP_1_port, A2 => A_EXP_1_port, ZN => 
                           n14384);
   U7530 : OAI21_X1 port map( B1 => n14407, B2 => n14385, A => n14384, ZN => 
                           n14406);
   U7531 : NAND2_X1 port map( A1 => n14505, A2 => n14473, ZN => n14386);
   U7532 : NAND2_X1 port map( A1 => n14406, A2 => n14386, ZN => n14388);
   U7533 : NAND2_X1 port map( A1 => B_EXP_2_port, A2 => A_EXP_2_port, ZN => 
                           n14387);
   U7534 : NAND2_X1 port map( A1 => n14388, A2 => n14387, ZN => n14404);
   U7535 : NAND2_X1 port map( A1 => n14504, A2 => n14472, ZN => n14389);
   U7536 : NAND2_X1 port map( A1 => n14404, A2 => n14389, ZN => n14391);
   U7537 : NAND2_X1 port map( A1 => B_EXP_3_port, A2 => A_EXP_3_port, ZN => 
                           n14390);
   U7538 : NAND2_X1 port map( A1 => n14391, A2 => n14390, ZN => n14410);
   U7539 : NAND2_X1 port map( A1 => n14506, A2 => n14475, ZN => n14393);
   U7540 : AND2_X1 port map( A1 => B_EXP_4_port, A2 => A_EXP_4_port, ZN => 
                           n14392);
   U7541 : AOI21_X1 port map( B1 => n14410, B2 => n14393, A => n14392, ZN => 
                           n14402);
   U7542 : NOR2_X1 port map( A1 => A_EXP_5_port, A2 => B_EXP_5_port, ZN => 
                           n14395);
   U7543 : NAND2_X1 port map( A1 => B_EXP_5_port, A2 => A_EXP_5_port, ZN => 
                           n14394);
   U7544 : OAI21_X1 port map( B1 => n14402, B2 => n14395, A => n14394, ZN => 
                           n14400);
   U7545 : NAND2_X1 port map( A1 => n14503, A2 => n14474, ZN => n14396);
   U7546 : AOI22_X1 port map( A1 => n14400, A2 => n14396, B1 => A_EXP_6_port, 
                           B2 => B_EXP_6_port, ZN => n14398);
   U7547 : XNOR2_X1 port map( A => B_EXP_7_port, B => A_EXP_7_port, ZN => 
                           n14397);
   U7548 : XNOR2_X1 port map( A => n14398, B => n14397, ZN => n374);
   U7549 : XNOR2_X1 port map( A => A_EXP_6_port, B => B_EXP_6_port, ZN => 
                           n14399);
   U7550 : XNOR2_X1 port map( A => n14400, B => n14399, ZN => 
                           I2_mw_I4sum_6_port);
   U7551 : XOR2_X1 port map( A => A_EXP_5_port, B => B_EXP_5_port, Z => n14401)
                           ;
   U7552 : XNOR2_X1 port map( A => n14402, B => n14401, ZN => 
                           I2_mw_I4sum_5_port);
   U7553 : XNOR2_X1 port map( A => A_EXP_3_port, B => B_EXP_3_port, ZN => 
                           n14403);
   U7554 : XNOR2_X1 port map( A => n14404, B => n14403, ZN => 
                           I2_mw_I4sum_3_port);
   U7555 : XNOR2_X1 port map( A => A_EXP_2_port, B => B_EXP_2_port, ZN => 
                           n14405);
   U7556 : XNOR2_X1 port map( A => n14406, B => n14405, ZN => 
                           I2_mw_I4sum_2_port);
   U7557 : XOR2_X1 port map( A => A_EXP_1_port, B => B_EXP_1_port, Z => n14408)
                           ;
   U7558 : XNOR2_X1 port map( A => n14408, B => n14407, ZN => 
                           I2_mw_I4sum_1_port);
   U7559 : XNOR2_X1 port map( A => A_EXP_4_port, B => B_EXP_4_port, ZN => 
                           n14409);
   U7560 : XNOR2_X1 port map( A => n14410, B => n14409, ZN => 
                           I2_mw_I4sum_4_port);
   U7561 : NOR2_X1 port map( A1 => n14416, A2 => n14493, ZN => n14418);
   U7562 : NAND2_X1 port map( A1 => n14418, A2 => n8376, ZN => n14411);
   U7563 : XNOR2_X1 port map( A => n14411, B => EXP_in_7_port, ZN => 
                           I3_EXP_out_7_port);
   U7564 : XNOR2_X1 port map( A => n14412, B => EXP_in_3_port, ZN => 
                           I3_EXP_out_3_port);
   U7565 : AND2_X1 port map( A1 => n14413, A2 => n2577, ZN => n14414);
   U7566 : NOR2_X1 port map( A1 => n14415, A2 => n14414, ZN => 
                           I3_EXP_out_1_port);
   U7567 : XNOR2_X1 port map( A => n14418, B => n14496, ZN => I3_EXP_out_6_port
                           );
   U7568 : AND2_X1 port map( A1 => n14416, A2 => n14493, ZN => n14417);
   U7569 : NOR2_X1 port map( A1 => n14418, A2 => n14417, ZN => 
                           I3_EXP_out_5_port);
   U7570 : NAND2_X1 port map( A1 => n14420, A2 => n14419, ZN => n14425);
   U7571 : NAND2_X1 port map( A1 => n14422, A2 => n14421, ZN => n14424);
   U7572 : MUX2_X1 port map( A => n14425, B => n14424, S => n14423, Z => n14427
                           );
   U7573 : NAND2_X1 port map( A1 => n14427, A2 => n14426, ZN => I1_isNaN_int);
   U7574 : INV_X1 port map( A => n14428, ZN => n14431);
   U7575 : AND2_X1 port map( A1 => n14446, A2 => n14429, ZN => n14430);
   U7576 : NAND3_X1 port map( A1 => n10847, A2 => n10812, A3 => n10846, ZN => 
                           n14922);
   U7577 : AND2_X1 port map( A1 => n14931, A2 => n14432, ZN => n14923);
   U7578 : XNOR2_X1 port map( A => n14926, B => EXP_out_round_2_port, ZN => 
                           n14433);
   U7579 : AND2_X1 port map( A1 => n14931, A2 => n14433, ZN => n14925);
   U7580 : OAI21_X1 port map( B1 => n14926, B2 => n14476, A => n14508, ZN => 
                           n14434);
   U7581 : INV_X1 port map( A => n14438, ZN => n14928);
   U7582 : XNOR2_X1 port map( A => n14438, B => n8379, ZN => n14437);
   U7583 : NAND2_X1 port map( A1 => n14438, A2 => n14498, ZN => n14439);
   U7584 : NAND2_X1 port map( A1 => n14439, A2 => n2579, ZN => n14440);
   U7585 : NAND3_X1 port map( A1 => n10812, A2 => n10833, A3 => n10832, ZN => 
                           n14930);
   U7586 : INV_X1 port map( A => FP_B(31), ZN => n14442);
   U7587 : XNOR2_X1 port map( A => n14442, B => FP_A(31), ZN => I1_SIGN_out_int
                           );
   U3762 : BUF_X1 port map( A => n11127, Z => n12837);
   U6485 : AOI21_X2 port map( B1 => n10694, B2 => n13026, A => n12995, ZN => 
                           n14079);
   U3969 : BUF_X1 port map( A => n14841, Z => n14121);
   U3944 : BUF_X2 port map( A => n11096, Z => n13979);
   U4040 : BUF_X1 port map( A => n14021, Z => n10940);
   U5184 : NOR2_X2 port map( A1 => n11899, A2 => n11898, ZN => n12915);
   U4130 : BUF_X2 port map( A => n11650, Z => n12805);
   I2_EXP_in_reg_6_inst : DFF_X1 port map( D => I2_EXP_in_tmp_6_port, CK => clk
                           , Q => n8376, QN => n14496);
   I2_EXP_in_reg_2_inst : DFF_X1 port map( D => I2_EXP_in_tmp_2_port, CK => clk
                           , Q => EXP_in_2_port, QN => n_1347);
   I2_EXP_in_tmp_reg_4_inst : DFF_X1 port map( D => I2_mw_I4sum_4_port, CK => 
                           clk, Q => n_1348, QN => n8323);
   R_1037 : DFFS_X1 port map( D => n14791, CK => clk, SN => n14950, Q => n14654
                           , QN => n_1349);
   R_1403 : DFFS_X1 port map( D => n14756, CK => clk, SN => n14949, Q => n14549
                           , QN => n_1350);
   R_1356 : DFFS_X1 port map( D => n14794, CK => clk, SN => n14948, Q => n14569
                           , QN => n_1351);
   R_1479 : SDFF_X1 port map( D => n12567, SI => n14947, SE => n12062, CK => 
                           clk, Q => n14020, QN => n_1352);
   U4166 : OR2_X2 port map( A1 => n11192, A2 => n11160, ZN => n11432);
   U4386 : AOI21_X2 port map( B1 => n13373, B2 => n14719, A => n14129, ZN => 
                           n11173);
   U3709 : BUF_X2 port map( A => n13221, Z => n14092);
   R_1284 : DFF_X2 port map( D => n14792, CK => clk, Q => n14598, QN => n_1353)
                           ;
   R_1487 : DFF_X1 port map( D => FP_B(14), CK => clk, Q => n14449, QN => 
                           n10869);
   R_1262 : DFF_X1 port map( D => n14606, CK => clk, Q => n14786, QN => n_1354)
                           ;
   U3685 : BUF_X1 port map( A => n12639, Z => n12142);
   U3590 : BUF_X1 port map( A => n11013, Z => n13347);
   U3600 : OR2_X1 port map( A1 => n10717, A2 => n10718, ZN => n13372);
   U3591 : BUF_X1 port map( A => n12125, Z => n11649);
   U4203 : NAND2_X1 port map( A1 => n10992, A2 => n10991, ZN => n12895);
   U3610 : AOI21_X1 port map( B1 => n11956, B2 => n13086, A => n11955, ZN => 
                           n13134);
   U3903 : OR3_X1 port map( A1 => n10928, A2 => n14675, A3 => n14674, ZN => 
                           n12490);
   U3907 : OR3_X1 port map( A1 => n10928, A2 => n14677, A3 => n14676, ZN => 
                           n12491);
   U4095 : OR3_X1 port map( A1 => n12488, A2 => n14665, A3 => n14664, ZN => 
                           n12492);
   U3582 : INV_X1 port map( A => n11823, ZN => n14964);
   U3583 : CLKBUF_X2 port map( A => n11127, Z => n13908);
   U3584 : XNOR2_X1 port map( A => n10855, B => n10854, ZN => 
                           intadd_47_SUM_3_port);
   U3589 : CLKBUF_X2 port map( A => n8339, Z => n13277);
   U3595 : BUF_X1 port map( A => n8353, Z => n11321);
   U3597 : CLKBUF_X1 port map( A => n8392, Z => n11965);
   U3599 : NOR2_X1 port map( A1 => n10598, A2 => n11324, ZN => n11504);
   U3602 : CLKBUF_X1 port map( A => n14780, Z => n12640);
   U3609 : CLKBUF_X1 port map( A => n14787, Z => n12018);
   U3612 : AND2_X1 port map( A1 => n10994, A2 => n10993, ZN => n12906);
   U3622 : CLKBUF_X1 port map( A => n8392, Z => n12743);
   U3626 : CLKBUF_X1 port map( A => n8392, Z => n13327);
   U3633 : BUF_X2 port map( A => n11237, Z => n12174);
   U3639 : NAND2_X1 port map( A1 => n11092, A2 => n11091, ZN => n11512);
   U3645 : XNOR2_X1 port map( A => n14648, B => n14649, ZN => n14954);
   U3654 : AND2_X1 port map( A1 => n11740, A2 => n11739, ZN => n11761);
   U3657 : BUF_X1 port map( A => n12783, Z => n13451);
   U3659 : CLKBUF_X2 port map( A => B_SIG_9_port, Z => n12764);
   U3662 : NAND2_X1 port map( A1 => n14941, A2 => n14940, ZN => n14953);
   U3666 : OR2_X1 port map( A1 => n12854, A2 => n12853, ZN => n12870);
   U3675 : CLKBUF_X2 port map( A => n8332, Z => n13234);
   U3679 : NAND2_X1 port map( A1 => n10600, A2 => n10599, ZN => n11634);
   U3686 : AND2_X1 port map( A1 => n12423, A2 => n10817, ZN => n12425);
   U3688 : XNOR2_X1 port map( A => intadd_47_SUM_3_port, B => n14954, ZN => 
                           intadd_46_SUM_4_port);
   U3729 : NOR2_X1 port map( A1 => n10627, A2 => n10625, ZN => n13294);
   U3755 : NOR2_X1 port map( A1 => n11890, A2 => n11889, ZN => n11989);
   U3770 : AND2_X1 port map( A1 => n12597, A2 => n12580, ZN => n13607);
   U3781 : NAND2_X1 port map( A1 => intadd_47_SUM_3_port, A2 => n14953, ZN => 
                           n14952);
   U3784 : BUF_X1 port map( A => n8332, Z => n12246);
   U3793 : NAND2_X1 port map( A1 => n14621, A2 => n10770, ZN => n14959);
   U3804 : OAI21_X1 port map( B1 => n14621, B2 => n10770, A => n14620, ZN => 
                           n14960);
   U3813 : NOR2_X1 port map( A1 => n12797, A2 => n12796, ZN => n13255);
   U3823 : NOR2_X1 port map( A1 => n12157, A2 => n12156, ZN => n12189);
   U3867 : NAND2_X1 port map( A1 => n14952, A2 => n14951, ZN => intadd_46_n1);
   U3875 : NAND2_X1 port map( A1 => n14960, A2 => n14959, ZN => n12388);
   U3884 : AOI22_X1 port map( A1 => n12399, A2 => n10784, B1 => n12398, B2 => 
                           n14647, ZN => n12607);
   U3885 : AND2_X1 port map( A1 => n13622, A2 => n13621, ZN => n11576);
   U3888 : AOI22_X1 port map( A1 => n13145, A2 => n13144, B1 => n13143, B2 => 
                           n13142, ZN => n14188);
   U3893 : NOR2_X1 port map( A1 => n14364, A2 => n10818, ZN => n13749);
   U3896 : XNOR2_X1 port map( A => n11791, B => n14964, ZN => n10906);
   U3906 : NAND2_X1 port map( A1 => n12386, A2 => n12385, ZN => n12597);
   U3908 : AND2_X1 port map( A1 => n12516, A2 => n14319, ZN => n12513);
   U3915 : CLKBUF_X1 port map( A => n12100, Z => n12265);
   U3916 : XNOR2_X1 port map( A => n13175, B => n14955, ZN => n13177);
   U3921 : CLKBUF_X1 port map( A => n14436, Z => n14438);
   U3940 : AND2_X1 port map( A1 => n14209, A2 => n14961, ZN => n10889);
   U3968 : OR3_X1 port map( A1 => n12100, A2 => n10789, A3 => n10758, ZN => 
                           n12342);
   U3977 : CLKBUF_X1 port map( A => n13731, Z => n13747);
   U3978 : OR3_X1 port map( A1 => n12488, A2 => n14665, A3 => n14664, ZN => 
                           n12489);
   U3985 : OR2_X1 port map( A1 => n14926, A2 => n12237, ZN => n14435);
   U4005 : NOR2_X1 port map( A1 => n2584, A2 => n12046, ZN => n14924);
   U4035 : CLKBUF_X1 port map( A => n12046, Z => n14446);
   U4042 : OR2_X1 port map( A1 => n10997, A2 => n10996, ZN => n12935);
   U4045 : INV_X1 port map( A => n14449, ZN => n14945);
   U4086 : XOR2_X1 port map( A => n11023, B => n11022, Z => n14946);
   U4087 : NAND2_X1 port map( A1 => n11839, A2 => n11838, ZN => n12033);
   n14947 <= '1';
   n14948 <= '1';
   n14949 <= '1';
   n14950 <= '1';
   U4126 : NAND2_X1 port map( A1 => n14648, A2 => n14649, ZN => n14951);
   U4156 : NAND2_X1 port map( A1 => n14957, A2 => n14956, ZN => n14955);
   U4159 : NAND2_X1 port map( A1 => n13172, A2 => n13173, ZN => n14956);
   U4167 : OAI21_X1 port map( B1 => n13173, B2 => n13172, A => n13174, ZN => 
                           n14957);
   U4175 : INV_X1 port map( A => n11512, ZN => n11510);
   U4176 : NAND3_X1 port map( A1 => n14943, A2 => n14944, A3 => n10787, ZN => 
                           n12100);
   U4177 : NAND4_X1 port map( A1 => n14958, A2 => n12415, A3 => n12409, A4 => 
                           n12412, ZN => n13688);
   U4209 : AND2_X1 port map( A1 => n12410, A2 => n12413, ZN => n14958);
   U4217 : OAI21_X1 port map( B1 => n11576, B2 => n13623, A => n13626, ZN => 
                           n11578);
   U4255 : NAND3_X1 port map( A1 => n12290, A2 => n12291, A3 => n14635, ZN => 
                           n12295);
   U4291 : OR2_X1 port map( A1 => n11729, A2 => n11730, ZN => n10960);
   U4350 : NAND2_X1 port map( A1 => n12033, A2 => n12034, ZN => n11843);
   U4606 : NAND3_X1 port map( A1 => n14206, A2 => n14205, A3 => n14962, ZN => 
                           n14961);
   U4740 : NAND2_X1 port map( A1 => n14963, A2 => n13550, ZN => n14962);
   U4741 : INV_X1 port map( A => n14207, ZN => n14963);
   U4742 : XNOR2_X1 port map( A => n13525, B => n10906, ZN => n10653);
   U4814 : NAND2_X1 port map( A1 => n11149, A2 => n13273, ZN => n11304);
   U4856 : XOR2_X1 port map( A => n10901, B => n13637, Z => n14965);

end SYN_pipeline;
