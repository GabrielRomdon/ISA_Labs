
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_FPmul is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_FPmul;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PackFP is

   port( SIGN : in std_logic;  EXP : in std_logic_vector (7 downto 0);  SIG : 
         in std_logic_vector (22 downto 0);  isNaN, isINF, isZ : in std_logic; 
         FP : out std_logic_vector (31 downto 0);  clk : in std_logic);

end PackFP;

architecture SYN_PackFP of PackFP is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal FP_22_port, FP_21_port, FP_20_port, FP_19_port, FP_18_port, 
      FP_17_port, FP_16_port, FP_15_port, FP_14_port, FP_13_port, FP_12_port, 
      FP_11_port, FP_10_port, FP_9_port, FP_8_port, FP_7_port, FP_6_port, 
      FP_5_port, FP_4_port, FP_3_port, FP_2_port, FP_1_port, FP_0_port, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n22, n23, n28, n29, n30, 
      FP_23_port, FP_24_port, FP_25_port, FP_26_port, FP_27_port, FP_28_port, 
      FP_29_port, FP_30_port, n39, n40, n47, n48, n67, n68, n70, n71, n72, n83,
      n84, n_1000, n_1001, n_1002, n_1003, n_1004 : std_logic;

begin
   FP <= ( SIGN, FP_30_port, FP_29_port, FP_28_port, FP_27_port, FP_26_port, 
      FP_25_port, FP_24_port, FP_23_port, FP_22_port, FP_21_port, FP_20_port, 
      FP_19_port, FP_18_port, FP_17_port, FP_16_port, FP_15_port, FP_14_port, 
      FP_13_port, FP_12_port, FP_11_port, FP_10_port, FP_9_port, FP_8_port, 
      FP_7_port, FP_6_port, FP_5_port, FP_4_port, FP_3_port, FP_2_port, 
      FP_1_port, FP_0_port );
   
   U20 : NAND2_X1 port map( A1 => SIG(22), A2 => n40, ZN => n23);
   U3 : NOR2_X1 port map( A1 => n71, A2 => n30, ZN => FP_9_port);
   U4 : NOR2_X1 port map( A1 => n72, A2 => n30, ZN => FP_8_port);
   U8 : INV_X1 port map( A => n22, ZN => FP_23_port);
   U10 : INV_X1 port map( A => n16, ZN => FP_28_port);
   U12 : INV_X1 port map( A => n19, ZN => FP_25_port);
   U13 : INV_X1 port map( A => n20, ZN => FP_24_port);
   U14 : INV_X1 port map( A => n18, ZN => FP_26_port);
   U15 : INV_X1 port map( A => n15, ZN => FP_29_port);
   U16 : INV_X1 port map( A => n17, ZN => FP_27_port);
   U17 : INV_X1 port map( A => n13, ZN => FP_30_port);
   U18 : INV_X1 port map( A => isZ, ZN => n39);
   U19 : AND2_X1 port map( A1 => n12, A2 => SIG(19), ZN => FP_19_port);
   U21 : AND2_X1 port map( A1 => n12, A2 => SIG(21), ZN => FP_21_port);
   U24 : AND2_X1 port map( A1 => n12, A2 => SIG(4), ZN => FP_4_port);
   U27 : AND2_X1 port map( A1 => n12, A2 => SIG(16), ZN => FP_16_port);
   U30 : AND2_X1 port map( A1 => n12, A2 => SIG(13), ZN => FP_13_port);
   U37 : AND2_X1 port map( A1 => n12, A2 => SIG(7), ZN => FP_7_port);
   U38 : INV_X1 port map( A => n12, ZN => n30);
   U39 : OAI21_X1 port map( B1 => n23, B2 => isZ, A => n67, ZN => FP_22_port);
   U40 : AOI21_X1 port map( B1 => EXP(7), B2 => n39, A => n14, ZN => n13);
   U41 : AOI21_X1 port map( B1 => EXP(6), B2 => n39, A => n14, ZN => n15);
   U42 : AOI21_X1 port map( B1 => EXP(5), B2 => n39, A => n14, ZN => n16);
   U43 : AOI21_X1 port map( B1 => EXP(4), B2 => n39, A => n14, ZN => n17);
   U44 : AOI21_X1 port map( B1 => EXP(3), B2 => n39, A => n14, ZN => n18);
   U45 : AOI21_X1 port map( B1 => EXP(2), B2 => n39, A => n14, ZN => n19);
   U46 : AOI21_X1 port map( B1 => EXP(1), B2 => n39, A => n14, ZN => n20);
   U47 : AOI21_X1 port map( B1 => EXP(0), B2 => n39, A => n14, ZN => n22);
   U48 : NOR2_X1 port map( A1 => isZ, A2 => n14, ZN => n28);
   U49 : NOR2_X1 port map( A1 => isZ, A2 => n14, ZN => n29);
   U29 : AND2_X1 port map( A1 => n28, A2 => SIG(14), ZN => FP_14_port);
   U28 : AND2_X1 port map( A1 => n29, A2 => SIG(15), ZN => FP_15_port);
   U26 : AND2_X1 port map( A1 => n28, A2 => SIG(17), ZN => FP_17_port);
   U25 : AND2_X1 port map( A1 => n29, A2 => SIG(18), ZN => FP_18_port);
   U22 : AND2_X1 port map( A1 => n29, A2 => SIG(20), ZN => FP_20_port);
   U31 : AND2_X1 port map( A1 => n29, A2 => SIG(12), ZN => FP_12_port);
   U11 : AND2_X1 port map( A1 => n28, A2 => SIG(2), ZN => FP_2_port);
   U33 : AND2_X1 port map( A1 => n29, A2 => SIG(10), ZN => FP_10_port);
   U7 : AND2_X1 port map( A1 => n28, A2 => SIG(5), ZN => FP_5_port);
   U23 : AND2_X1 port map( A1 => n28, A2 => SIG(1), ZN => FP_1_port);
   U9 : AND2_X1 port map( A1 => n29, A2 => SIG(3), ZN => FP_3_port);
   U6 : AND2_X1 port map( A1 => n29, A2 => SIG(6), ZN => FP_6_port);
   U32 : NOR2_X1 port map( A1 => isZ, A2 => n14, ZN => n12);
   U34 : AND2_X1 port map( A1 => n28, A2 => SIG(0), ZN => FP_0_port);
   U35 : AND2_X1 port map( A1 => n28, A2 => SIG(11), ZN => FP_11_port);
   U51 : INV_X1 port map( A => SIG(8), ZN => n47);
   U52 : INV_X1 port map( A => SIG(9), ZN => n48);
   U5 : INV_X1 port map( A => isINF, ZN => n40);
   U36 : OR2_X1 port map( A1 => isINF, A2 => n84, ZN => n14);
   MY_CLK_r_REG1031_S3 : DFF_X1 port map( D => n70, CK => clk, Q => n_1000, QN 
                           => n83);
   MY_CLK_r_REG1033_S5 : DFF_X1 port map( D => n68, CK => clk, Q => n67, QN => 
                           n84);
   MY_CLK_r_REG1049_S5 : DFF_X1 port map( D => n48, CK => clk, Q => n71, QN => 
                           n_1001);
   MY_CLK_r_REG1046_S5 : DFF_X1 port map( D => n47, CK => clk, Q => n72, QN => 
                           n_1002);
   MY_CLK_r_REG1032_S4 : DFF_X1 port map( D => n83, CK => clk, Q => n68, QN => 
                           n_1003);
   MY_CLK_r_REG1030_S2 : DFF_X1 port map( D => isNaN, CK => clk, Q => n70, QN 
                           => n_1004);

end SYN_PackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPnormalize_SIG_width28_1 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
         std_logic);

end FPnormalize_SIG_width28_1;

architecture SYN_FPnormalize of FPnormalize_SIG_width28_1 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n21, n22, n23, n24, n25, n153, n167, n168, n169, n171, n172, n173, 
      n174, n255, n256, n257, n258, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n363, n364, n365, n366, n367, n_1012, n_1013, n_1014, 
      n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028 : std_logic;

begin
   
   U34 : MUX2_X1 port map( A => n295, B => SIG_in(9), S => n255, Z => 
                           SIG_out(9));
   U35 : MUX2_X1 port map( A => SIG_in(9), B => SIG_in(8), S => n255, Z => 
                           SIG_out(8));
   U36 : MUX2_X1 port map( A => SIG_in(8), B => SIG_in(7), S => n255, Z => 
                           SIG_out(7));
   U37 : MUX2_X1 port map( A => SIG_in(7), B => SIG_in(6), S => n255, Z => 
                           SIG_out(6));
   U38 : MUX2_X1 port map( A => SIG_in(6), B => SIG_in(5), S => n255, Z => 
                           SIG_out(5));
   U39 : MUX2_X1 port map( A => SIG_in(5), B => SIG_in(4), S => n255, Z => 
                           SIG_out(4));
   U40 : MUX2_X1 port map( A => SIG_in(4), B => SIG_in(3), S => n255, Z => 
                           SIG_out(3));
   U41 : MUX2_X1 port map( A => SIG_in(26), B => SIG_in(25), S => n255, Z => 
                           SIG_out(25));
   U42 : MUX2_X1 port map( A => SIG_in(25), B => SIG_in(24), S => n255, Z => 
                           SIG_out(24));
   U43 : MUX2_X1 port map( A => SIG_in(24), B => SIG_in(23), S => n255, Z => 
                           SIG_out(23));
   U44 : MUX2_X1 port map( A => SIG_in(23), B => SIG_in(22), S => n255, Z => 
                           SIG_out(22));
   U45 : MUX2_X1 port map( A => SIG_in(22), B => SIG_in(21), S => n255, Z => 
                           SIG_out(21));
   U46 : MUX2_X1 port map( A => SIG_in(21), B => SIG_in(20), S => n255, Z => 
                           SIG_out(20));
   U47 : MUX2_X1 port map( A => SIG_in(20), B => SIG_in(19), S => n255, Z => 
                           SIG_out(19));
   U48 : MUX2_X1 port map( A => SIG_in(19), B => SIG_in(18), S => n255, Z => 
                           SIG_out(18));
   U49 : MUX2_X1 port map( A => SIG_in(18), B => SIG_in(17), S => n255, Z => 
                           SIG_out(17));
   U50 : MUX2_X1 port map( A => SIG_in(17), B => SIG_in(16), S => n255, Z => 
                           SIG_out(16));
   U51 : MUX2_X1 port map( A => SIG_in(16), B => SIG_in(15), S => n255, Z => 
                           SIG_out(15));
   U52 : MUX2_X1 port map( A => SIG_in(15), B => n299, S => n255, Z => 
                           SIG_out(14));
   U53 : MUX2_X1 port map( A => n299, B => n298, S => n255, Z => SIG_out(13));
   U54 : MUX2_X1 port map( A => n298, B => n297, S => n255, Z => SIG_out(12));
   U55 : MUX2_X1 port map( A => n297, B => n296, S => n255, Z => SIG_out(11));
   U56 : MUX2_X1 port map( A => n296, B => n295, S => n255, Z => SIG_out(10));
   U57 : XOR2_X1 port map( A => n286, B => n258, Z => EXP_out(4));
   U58 : XOR2_X1 port map( A => n300, B => n283, Z => EXP_out(3));
   U59 : XOR2_X1 port map( A => n302, B => n24, Z => EXP_out(2));
   U3 : OR2_X1 port map( A1 => SIG_in(27), A2 => SIG_in(26), ZN => SIG_out(26))
                           ;
   U13 : NOR2_X1 port map( A1 => n365, A2 => n255, ZN => n25);
   U12 : XNOR2_X1 port map( A => n303, B => n25, ZN => EXP_out(1));
   U14 : AOI22_X1 port map( A1 => SIG_in(27), A2 => n294, B1 => n365, B2 => 
                           n255, ZN => EXP_out(0));
   U6 : XNOR2_X1 port map( A => n290, B => n22, ZN => EXP_out(6));
   U8 : XNOR2_X1 port map( A => n292, B => n23, ZN => EXP_out(5));
   U30 : NOR2_X1 port map( A1 => n286, A2 => n258, ZN => n23);
   U31 : XNOR2_X1 port map( A => n288, B => n21, ZN => EXP_out(7));
   U32 : NOR3_X1 port map( A1 => n286, A2 => n292, A3 => n258, ZN => n22);
   U10 : OR2_X1 port map( A1 => n302, A2 => n24, ZN => n153);
   U77 : INV_X1 port map( A => EXP_in(1), ZN => n167);
   U78 : INV_X1 port map( A => EXP_in(2), ZN => n168);
   U79 : INV_X1 port map( A => EXP_in(3), ZN => n169);
   U2 : OR3_X1 port map( A1 => n303, A2 => n365, A3 => n255, ZN => n24);
   U7 : NOR2_X1 port map( A1 => n258, A2 => n282, ZN => n21);
   U9 : NAND2_X1 port map( A1 => n285, A2 => n284, ZN => n258);
   U15 : NAND3_X1 port map( A1 => n363, A2 => n364, A3 => n367, ZN => n256);
   MY_CLK_r_REG1085_S4 : DFF_X1 port map( D => n169, CK => clk, Q => n301, QN 
                           => n366);
   MY_CLK_r_REG1105_S4 : DFF_X1 port map( D => EXP_in(0), CK => clk, Q => n294,
                           QN => n365);
   MY_CLK_r_REG1095_S4 : DFF_X1 port map( D => n171, CK => clk, Q => n293, QN 
                           => n367);
   MY_CLK_r_REG1093_S4 : DFF_X1 port map( D => n172, CK => clk, Q => n291, QN 
                           => n364);
   MY_CLK_r_REG1088_S4 : DFF_X1 port map( D => n174, CK => clk, Q => n287, QN 
                           => n363);
   U21 : INV_X1 port map( A => n153, ZN => n257);
   U23 : INV_X1 port map( A => EXP_in(4), ZN => n174);
   U24 : INV_X1 port map( A => EXP_in(7), ZN => n173);
   U25 : INV_X1 port map( A => EXP_in(6), ZN => n172);
   U27 : INV_X1 port map( A => EXP_in(5), ZN => n171);
   U4 : INV_X2 port map( A => SIG_in(27), ZN => n255);
   MY_CLK_r_REG1112_S4 : DFF_X1 port map( D => n167, CK => clk, Q => n303, QN 
                           => n_1012);
   MY_CLK_r_REG1096_S5 : DFF_X1 port map( D => n293, CK => clk, Q => n292, QN 
                           => n_1013);
   MY_CLK_r_REG1094_S5 : DFF_X1 port map( D => n291, CK => clk, Q => n290, QN 
                           => n_1014);
   MY_CLK_r_REG1092_S5 : DFF_X1 port map( D => n289, CK => clk, Q => n288, QN 
                           => n_1015);
   MY_CLK_r_REG1091_S4 : DFF_X1 port map( D => n173, CK => clk, Q => n289, QN 
                           => n_1016);
   MY_CLK_r_REG1090_S5 : DFF_X1 port map( D => n256, CK => clk, Q => n282, QN 
                           => n_1017);
   MY_CLK_r_REG1089_S5 : DFF_X1 port map( D => n287, CK => clk, Q => n286, QN 
                           => n_1018);
   MY_CLK_r_REG1087_S5 : DFF_X1 port map( D => n366, CK => clk, Q => n284, QN 
                           => n_1019);
   MY_CLK_r_REG1086_S5 : DFF_X1 port map( D => n301, CK => clk, Q => n300, QN 
                           => n_1020);
   MY_CLK_r_REG1084_S4 : DFF_X1 port map( D => n168, CK => clk, Q => n302, QN 
                           => n_1021);
   MY_CLK_r_REG1080_S4 : DFF_X1 port map( D => SIG_in(10), CK => clk, Q => n295
                           , QN => n_1022);
   MY_CLK_r_REG1069_S5 : DFF_X1 port map( D => n257, CK => clk, Q => n285, QN 
                           => n_1023);
   MY_CLK_r_REG1068_S5 : DFF_X1 port map( D => n153, CK => clk, Q => n283, QN 
                           => n_1024);
   MY_CLK_r_REG1052_S4 : DFF_X1 port map( D => SIG_in(14), CK => clk, Q => n299
                           , QN => n_1025);
   MY_CLK_r_REG1050_S4 : DFF_X1 port map( D => SIG_in(13), CK => clk, Q => n298
                           , QN => n_1026);
   MY_CLK_r_REG1048_S4 : DFF_X1 port map( D => SIG_in(12), CK => clk, Q => n297
                           , QN => n_1027);
   MY_CLK_r_REG1044_S4 : DFF_X1 port map( D => SIG_in(11), CK => clk, Q => n296
                           , QN => n_1028);

end SYN_FPnormalize;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPround_SIG_width28 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
         std_logic);

end FPround_SIG_width28;

architecture SYN_FPround of FPround_SIG_width28 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal N5, N6, N7, N8, N10, N11, N12, N13, N14, N15, N16, N18, N19, n122, 
      n36, n48, n53, add_45_n24, add_45_n23, add_45_n19, add_45_n15, add_45_n14
      , add_45_carry_3_port, add_45_carry_5_port, add_45_carry_6_port, 
      add_45_carry_7_port, add_45_carry_10_port, add_45_carry_11_port, 
      add_45_carry_12_port, add_45_carry_14_port, add_45_carry_15_port, 
      add_45_carry_18_port, add_45_carry_21_port, add_45_carry_22_port, 
      add_45_carry_23_port, n177, n179, n188, n194, n195, n196, n197, n198, 
      n199, n200, n201, n203, n204, n205, n212, n213, n229, n230, n339, n340, 
      n349, n350, n354, n355, n356, n357, n360, n362, n363, n364, n365, n366, 
      n368, n369, n370, n372, n374, n401, n402, n403, n404, n405, n406, n407, 
      n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, 
      n420, n422, n423, n424, n425, n455, n456, n457, n458, n459, n460, n461, 
      n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, 
      n474, n476, n477, n480, n481, n482, n484, n485, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041 : std_logic;

begin
   EXP_out <= ( EXP_in(7), EXP_in(6), EXP_in(5), EXP_in(4), EXP_in(3), 
      EXP_in(2), EXP_in(1), EXP_in(0) );
   
   add_45_U2 : AND2_X1 port map( A1 => n403, A2 => n415, ZN => n230);
   add_45_U11 : AND2_X1 port map( A1 => n230, A2 => n416, ZN => add_45_n23);
   add_45_U21 : XNOR2_X1 port map( A => n213, B => add_45_n14, ZN => N10);
   add_45_U30 : XNOR2_X1 port map( A => add_45_carry_14_port, B => n458, ZN => 
                           N16);
   add_45_U16 : XNOR2_X1 port map( A => n403, B => n459, ZN => n229);
   add_45_U19 : XNOR2_X1 port map( A => add_45_n23, B => n466, ZN => N19);
   add_45_U1_1_3 : HA_X1 port map( A => n409, B => n188, CO => add_45_n19, S =>
                           N5);
   add_45_U1_1_4 : HA_X1 port map( A => add_45_n19, B => n410, CO => 
                           add_45_carry_5_port, S => N6);
   add_45_U1_1_5 : HA_X1 port map( A => add_45_carry_5_port, B => n411, CO => 
                           add_45_carry_6_port, S => N7);
   add_45_U1_1_6 : HA_X1 port map( A => add_45_carry_6_port, B => n412, CO => 
                           n_1035, S => N8);
   U5 : NAND2_X1 port map( A1 => SIG_in(9), A2 => SIG_in(7), ZN => n177);
   U10 : AND2_X1 port map( A1 => n407, A2 => n464, ZN => add_45_n24);
   U13 : AND2_X1 port map( A1 => add_45_n24, A2 => n408, ZN => n188);
   U25 : AOI22_X1 port map( A1 => n405, A2 => n464, B1 => n404, B2 => n425, ZN 
                           => SIG_out(3));
   U26 : AOI22_X1 port map( A1 => SIG_in(2), A2 => n349, B1 => n122, B2 => n36,
                           ZN => SIG_out(10));
   U27 : AOI22_X1 port map( A1 => n406, A2 => n340, B1 => n404, B2 => n455, ZN 
                           => SIG_out(4));
   U28 : AOI22_X1 port map( A1 => n406, A2 => n48, B1 => n404, B2 => n472, ZN 
                           => SIG_out(6));
   U29 : AOI22_X1 port map( A1 => n405, A2 => n339, B1 => n404, B2 => n469, ZN 
                           => SIG_out(5));
   U30 : OAI21_X1 port map( B1 => n406, B2 => n456, A => n194, ZN => SIG_out(7)
                           );
   U31 : NAND2_X1 port map( A1 => N6, A2 => n405, ZN => n194);
   U32 : OAI21_X1 port map( B1 => n406, B2 => n468, A => n195, ZN => SIG_out(8)
                           );
   U33 : NAND2_X1 port map( A1 => N7, A2 => n405, ZN => n195);
   U34 : OAI21_X1 port map( B1 => SIG_in(2), B2 => n368, A => n197, ZN => 
                           SIG_out(12));
   U35 : NAND2_X1 port map( A1 => N11, A2 => SIG_in(2), ZN => n197);
   U36 : OAI21_X1 port map( B1 => SIG_in(2), B2 => n362, A => n198, ZN => 
                           SIG_out(13));
   U37 : NAND2_X1 port map( A1 => N12, A2 => SIG_in(2), ZN => n198);
   U38 : OAI21_X1 port map( B1 => n406, B2 => n457, A => n196, ZN => SIG_out(9)
                           );
   U39 : NAND2_X1 port map( A1 => N8, A2 => n406, ZN => n196);
   U40 : OAI21_X1 port map( B1 => SIG_in(2), B2 => n363, A => n199, ZN => 
                           SIG_out(14));
   U41 : NAND2_X1 port map( A1 => N13, A2 => SIG_in(2), ZN => n199);
   U42 : OAI21_X1 port map( B1 => n405, B2 => n424, A => n200, ZN => 
                           SIG_out(15));
   U43 : NAND2_X1 port map( A1 => n402, A2 => n406, ZN => n200);
   U44 : OAI21_X1 port map( B1 => n405, B2 => n467, A => n201, ZN => 
                           SIG_out(16));
   U45 : NAND2_X1 port map( A1 => N15, A2 => n405, ZN => n201);
   U46 : OAI22_X1 port map( A1 => n356, A2 => n471, B1 => n470, B2 => n473, ZN 
                           => SIG_out(25));
   U47 : OAI22_X1 port map( A1 => n354, A2 => n471, B1 => n470, B2 => n463, ZN 
                           => SIG_out(23));
   U48 : OAI22_X1 port map( A1 => n355, A2 => n471, B1 => n470, B2 => n477, ZN 
                           => SIG_out(24));
   U49 : OAI22_X1 port map( A1 => n471, A2 => n350, B1 => n470, B2 => n461, ZN 
                           => SIG_out(21));
   U50 : OAI22_X1 port map( A1 => n212, A2 => n471, B1 => n470, B2 => n462, ZN 
                           => SIG_out(22));
   U53 : OAI21_X1 port map( B1 => n406, B2 => n459, A => n203, ZN => 
                           SIG_out(18));
   U54 : NAND2_X1 port map( A1 => n229, A2 => n406, ZN => n203);
   U55 : OAI22_X1 port map( A1 => n357, A2 => n471, B1 => n465, B2 => n470, ZN 
                           => SIG_out(26));
   U56 : OAI21_X1 port map( B1 => n466, B2 => n406, A => n205, ZN => 
                           SIG_out(20));
   U57 : NAND2_X1 port map( A1 => N19, A2 => n406, ZN => n205);
   U58 : OAI21_X1 port map( B1 => n406, B2 => n460, A => n204, ZN => 
                           SIG_out(19));
   U59 : NAND2_X1 port map( A1 => N18, A2 => n406, ZN => n204);
   U60 : MUX2_X1 port map( A => N10, B => SIG_in(11), S => n122, Z => 
                           SIG_out(11));
   U3 : XOR2_X1 port map( A => n462, B => add_45_n15, Z => n212);
   U4 : AND3_X1 port map( A1 => SIG_in(5), A2 => SIG_in(3), A3 => SIG_in(4), ZN
                           => add_45_carry_3_port);
   U76 : INV_X1 port map( A => SIG_in(10), ZN => n36);
   U78 : INV_X1 port map( A => N5, ZN => n48);
   U89 : INV_X1 port map( A => SIG_in(11), ZN => n213);
   U92 : INV_X1 port map( A => SIG_in(3), ZN => n53);
   add_45_U32 : AND2_X1 port map( A1 => add_45_carry_18_port, A2 => n418, ZN =>
                           add_45_n15);
   U8 : AND2_X1 port map( A1 => add_45_carry_11_port, A2 => SIG_in(14), ZN => 
                           add_45_carry_12_port);
   U14 : AND2_X1 port map( A1 => add_45_carry_22_port, A2 => n422, ZN => 
                           add_45_carry_23_port);
   U17 : AND2_X1 port map( A1 => add_45_carry_7_port, A2 => SIG_in(10), ZN => 
                           add_45_n14);
   U19 : NOR2_X1 port map( A1 => n179, A2 => n177, ZN => add_45_carry_7_port);
   U20 : NOR2_X1 port map( A1 => n366, A2 => n463, ZN => add_45_carry_21_port);
   U21 : NAND2_X1 port map( A1 => add_45_n15, A2 => n419, ZN => n366);
   U22 : AND2_X1 port map( A1 => n423, A2 => n406, ZN => n364);
   U51 : XOR2_X1 port map( A => add_45_n24, B => n469, Z => n339);
   U52 : XNOR2_X1 port map( A => n407, B => n464, ZN => n340);
   U62 : XOR2_X1 port map( A => add_45_carry_7_port, B => n36, Z => n349);
   U63 : XOR2_X1 port map( A => add_45_carry_18_port, B => n461, Z => n350);
   U64 : XOR2_X1 port map( A => n366, B => n420, Z => n354);
   U65 : XOR2_X1 port map( A => add_45_carry_21_port, B => n477, Z => n355);
   U66 : XOR2_X1 port map( A => add_45_carry_22_port, B => n473, Z => n356);
   U68 : XOR2_X1 port map( A => add_45_carry_23_port, B => n465, Z => n357);
   U77 : AND2_X1 port map( A1 => SIG_in(15), A2 => SIG_in(14), ZN => n360);
   U80 : AND2_X1 port map( A1 => n401, A2 => n413, ZN => add_45_carry_14_port);
   U81 : XNOR2_X1 port map( A => add_45_carry_12_port, B => n365, ZN => N14);
   U82 : XNOR2_X1 port map( A => n401, B => n467, ZN => N15);
   U85 : XNOR2_X1 port map( A => add_45_carry_10_port, B => n362, ZN => N12);
   U86 : INV_X1 port map( A => SIG_in(13), ZN => n362);
   U87 : NAND2_X1 port map( A1 => add_45_n14, A2 => SIG_in(11), ZN => n369);
   U88 : XNOR2_X1 port map( A => add_45_carry_11_port, B => n363, ZN => N13);
   U90 : INV_X1 port map( A => SIG_in(14), ZN => n363);
   U91 : INV_X1 port map( A => SIG_in(15), ZN => n365);
   U93 : XNOR2_X1 port map( A => n460, B => n230, ZN => N18);
   U95 : INV_X1 port map( A => SIG_in(12), ZN => n368);
   U96 : XNOR2_X1 port map( A => n369, B => SIG_in(12), ZN => N11);
   U97 : NAND2_X1 port map( A1 => n372, A2 => n370, ZN => SIG_out(17));
   U98 : NAND2_X1 port map( A1 => n404, A2 => n414, ZN => n370);
   U99 : NAND2_X1 port map( A1 => N16, A2 => n406, ZN => n372);
   U12 : AND3_X1 port map( A1 => add_45_carry_10_port, A2 => n360, A3 => 
                           SIG_in(13), ZN => n374);
   U15 : INV_X1 port map( A => SIG_in(2), ZN => n122);
   U18 : NAND3_X1 port map( A1 => add_45_carry_3_port, A2 => SIG_in(6), A3 => 
                           SIG_in(8), ZN => n179);
   MY_CLK_r_REG1081_S4 : DFF_X1 port map( D => n53, CK => clk, Q => n425, QN =>
                           n464);
   MY_CLK_r_REG1100_S4 : DFF_X1 port map( D => SIG_in(26), CK => clk, Q => n423
                           , QN => n465);
   MY_CLK_r_REG1113_S4 : DFF_X1 port map( D => SIG_in(25), CK => clk, Q => n422
                           , QN => n473);
   MY_CLK_r_REG1111_S4 : DFF_X1 port map( D => SIG_in(24), CK => clk, Q => 
                           n_1036, QN => n477);
   MY_CLK_r_REG1115_S4 : DFF_X1 port map( D => SIG_in(23), CK => clk, Q => n420
                           , QN => n463);
   MY_CLK_r_REG1103_S4 : DFF_X1 port map( D => SIG_in(22), CK => clk, Q => n419
                           , QN => n462);
   MY_CLK_r_REG1101_S4 : DFF_X1 port map( D => SIG_in(21), CK => clk, Q => n418
                           , QN => n461);
   MY_CLK_r_REG1114_S4 : DFF_X1 port map( D => SIG_in(20), CK => clk, Q => n417
                           , QN => n466);
   MY_CLK_r_REG1104_S4 : DFF_X1 port map( D => SIG_in(19), CK => clk, Q => n416
                           , QN => n460);
   MY_CLK_r_REG1107_S4 : DFF_X1 port map( D => SIG_in(18), CK => clk, Q => n415
                           , QN => n459);
   MY_CLK_r_REG1102_S4 : DFF_X1 port map( D => SIG_in(17), CK => clk, Q => n414
                           , QN => n458);
   MY_CLK_r_REG1116_S4 : DFF_X1 port map( D => SIG_in(16), CK => clk, Q => n413
                           , QN => n467);
   MY_CLK_r_REG1097_S4 : DFF_X1 port map( D => SIG_in(9), CK => clk, Q => n412,
                           QN => n457);
   MY_CLK_r_REG1098_S4 : DFF_X1 port map( D => SIG_in(8), CK => clk, Q => n411,
                           QN => n468);
   MY_CLK_r_REG1083_S4 : DFF_X1 port map( D => SIG_in(7), CK => clk, Q => n410,
                           QN => n456);
   MY_CLK_r_REG1099_S4 : DFF_X1 port map( D => SIG_in(6), CK => clk, Q => n409,
                           QN => n472);
   MY_CLK_r_REG1082_S4 : DFF_X1 port map( D => SIG_in(5), CK => clk, Q => n408,
                           QN => n469);
   MY_CLK_r_REG1043_S4 : DFF_X1 port map( D => SIG_in(4), CK => clk, Q => n407,
                           QN => n455);
   MY_CLK_r_REG1108_S4 : DFF_X1 port map( D => SIG_in(2), CK => clk, Q => n406,
                           QN => n471);
   MY_CLK_r_REG1109_S4 : DFF_X1 port map( D => n122, CK => clk, Q => n404, QN 
                           => n470);
   U6 : NOR2_X1 port map( A1 => n369, A2 => n368, ZN => add_45_carry_10_port);
   U7 : NOR2_X1 port map( A1 => n474, A2 => n369, ZN => add_45_carry_11_port);
   U9 : NAND2_X1 port map( A1 => SIG_in(13), A2 => SIG_in(12), ZN => n474);
   U61 : OR2_X1 port map( A1 => n477, A2 => n463, ZN => n476);
   U67 : NOR2_X1 port map( A1 => n482, A2 => n481, ZN => n480);
   U69 : AND2_X1 port map( A1 => n374, A2 => n480, ZN => add_45_carry_15_port);
   U70 : INV_X1 port map( A => SIG_in(17), ZN => n481);
   U71 : INV_X1 port map( A => SIG_in(16), ZN => n482);
   U11 : NOR2_X1 port map( A1 => n476, A2 => n462, ZN => n484);
   U16 : AND2_X1 port map( A1 => n417, A2 => n416, ZN => n485);
   U23 : AND2_X1 port map( A1 => n230, A2 => n485, ZN => add_45_carry_18_port);
   U24 : AND2_X1 port map( A1 => add_45_n15, A2 => n484, ZN => 
                           add_45_carry_22_port);
   U72 : AND2_X1 port map( A1 => add_45_carry_23_port, A2 => n364, ZN => 
                           SIG_out(27));
   MY_CLK_r_REG1110_S4 : DFF_X1 port map( D => SIG_in(2), CK => clk, Q => n405,
                           QN => n_1037);
   MY_CLK_r_REG1106_S4 : DFF_X1 port map( D => n365, CK => clk, Q => n424, QN 
                           => n_1038);
   MY_CLK_r_REG1057_S4 : DFF_X1 port map( D => add_45_carry_15_port, CK => clk,
                           Q => n403, QN => n_1039);
   MY_CLK_r_REG1056_S4 : DFF_X1 port map( D => n374, CK => clk, Q => n401, QN 
                           => n_1040);
   MY_CLK_r_REG1054_S4 : DFF_X1 port map( D => N14, CK => clk, Q => n402, QN =>
                           n_1041);

end SYN_FPround;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPnormalize_SIG_width28_0 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
         std_logic);

end FPnormalize_SIG_width28_0;

architecture SYN_FPnormalize of FPnormalize_SIG_width28_0 is

   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n52, n61, n63, n162, n167, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n237, n238, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087 : std_logic;

begin
   
   U10 : XNOR2_X1 port map( A => n230, B => n4, ZN => EXP_out(3));
   U19 : MUX2_X1 port map( A => n244, B => n245, S => n345, Z => SIG_out(9));
   U20 : MUX2_X1 port map( A => n243, B => n244, S => n345, Z => SIG_out(8));
   U21 : MUX2_X1 port map( A => n242, B => n243, S => n345, Z => SIG_out(7));
   U27 : MUX2_X1 port map( A => n256, B => SIG_in(26), S => n52, Z => 
                           SIG_out(25));
   U28 : MUX2_X1 port map( A => n255, B => n256, S => n52, Z => SIG_out(24));
   U29 : MUX2_X1 port map( A => n254, B => n255, S => n52, Z => SIG_out(23));
   U30 : MUX2_X1 port map( A => SIG_in(22), B => n254, S => n52, Z => 
                           SIG_out(22));
   U31 : MUX2_X1 port map( A => SIG_in(21), B => SIG_in(22), S => n52, Z => 
                           SIG_out(21));
   U32 : MUX2_X1 port map( A => SIG_in(20), B => SIG_in(21), S => n52, Z => 
                           SIG_out(20));
   U33 : MUX2_X1 port map( A => SIG_in(19), B => SIG_in(20), S => n52, Z => 
                           SIG_out(19));
   U34 : MUX2_X1 port map( A => n253, B => SIG_in(19), S => n52, Z => 
                           SIG_out(18));
   U35 : MUX2_X1 port map( A => n252, B => n253, S => n52, Z => SIG_out(17));
   U36 : MUX2_X1 port map( A => n251, B => n252, S => n52, Z => SIG_out(16));
   U37 : MUX2_X1 port map( A => n250, B => n251, S => n52, Z => SIG_out(15));
   U38 : MUX2_X1 port map( A => n249, B => n250, S => n52, Z => SIG_out(14));
   U39 : MUX2_X1 port map( A => n248, B => n249, S => n52, Z => SIG_out(13));
   U40 : MUX2_X1 port map( A => n247, B => n248, S => n52, Z => SIG_out(12));
   U41 : MUX2_X1 port map( A => n246, B => n247, S => n52, Z => SIG_out(11));
   U42 : MUX2_X1 port map( A => n245, B => n246, S => n52, Z => SIG_out(10));
   U43 : XOR2_X1 port map( A => n219, B => n162, Z => EXP_out(4));
   U44 : XOR2_X1 port map( A => n8, B => n227, Z => EXP_out(2));
   U13 : XNOR2_X1 port map( A => n224, B => n9, ZN => EXP_out(1));
   U5 : NOR4_X1 port map( A1 => n215, A2 => n219, A3 => n217, A4 => n162, ZN =>
                           n5);
   U4 : XNOR2_X1 port map( A => n213, B => n5, ZN => EXP_out(7));
   U7 : NOR3_X1 port map( A1 => n219, A2 => n217, A3 => n162, ZN => n6);
   U6 : XNOR2_X1 port map( A => n215, B => n6, ZN => EXP_out(6));
   U9 : NOR2_X1 port map( A1 => n219, A2 => n162, ZN => n7);
   U8 : XNOR2_X1 port map( A => n217, B => n7, ZN => EXP_out(5));
   U3 : OR2_X1 port map( A1 => n52, A2 => SIG_in(26), ZN => SIG_out(26));
   U48 : AOI22_X1 port map( A1 => n52, A2 => n221, B1 => n339, B2 => n167, ZN 
                           => EXP_out(0));
   U49 : NAND2_X1 port map( A1 => n52, A2 => n221, ZN => n9);
   U50 : OAI21_X1 port map( B1 => n343, B2 => n345, A => n63, ZN => SIG_out(4))
                           ;
   U51 : OAI21_X1 port map( B1 => n337, B2 => n345, A => n61, ZN => SIG_out(3))
                           ;
   U52 : NAND2_X1 port map( A1 => SIG_in(27), A2 => n240, ZN => n63);
   U54 : MUX2_X1 port map( A => n240, B => n241, S => n345, Z => SIG_out(5));
   U12 : AND3_X1 port map( A1 => n345, A2 => n221, A3 => n224, ZN => n8);
   U11 : NAND2_X1 port map( A1 => n8, A2 => n227, ZN => n4);
   U22 : MUX2_X1 port map( A => n241, B => n242, S => n345, Z => SIG_out(6));
   U16 : MUX2_X1 port map( A => n237, B => n238, S => n52, Z => SIG_out(2));
   U18 : OR2_X1 port map( A1 => n167, A2 => n343, ZN => n61);
   MY_CLK_r_REG1118_S3 : DFF_X1 port map( D => SIG_in(25), CK => clk, Q => n256
                           , QN => n_1047);
   MY_CLK_r_REG1119_S3 : DFF_X1 port map( D => SIG_in(24), CK => clk, Q => n255
                           , QN => n_1048);
   MY_CLK_r_REG1120_S3 : DFF_X1 port map( D => SIG_in(23), CK => clk, Q => n254
                           , QN => n_1049);
   MY_CLK_r_REG1123_S3 : DFF_X1 port map( D => SIG_in(18), CK => clk, Q => n253
                           , QN => n_1050);
   MY_CLK_r_REG1128_S3 : DFF_X1 port map( D => SIG_in(17), CK => clk, Q => n252
                           , QN => n_1051);
   MY_CLK_r_REG1127_S3 : DFF_X1 port map( D => SIG_in(16), CK => clk, Q => n251
                           , QN => n_1052);
   MY_CLK_r_REG1130_S3 : DFF_X1 port map( D => SIG_in(15), CK => clk, Q => n250
                           , QN => n_1053);
   MY_CLK_r_REG1129_S3 : DFF_X1 port map( D => SIG_in(14), CK => clk, Q => n249
                           , QN => n_1054);
   MY_CLK_r_REG1134_S3 : DFF_X1 port map( D => SIG_in(13), CK => clk, Q => n248
                           , QN => n_1055);
   MY_CLK_r_REG1133_S3 : DFF_X1 port map( D => SIG_in(12), CK => clk, Q => n247
                           , QN => n_1056);
   MY_CLK_r_REG1131_S3 : DFF_X1 port map( D => SIG_in(11), CK => clk, Q => n246
                           , QN => n_1057);
   MY_CLK_r_REG1132_S3 : DFF_X1 port map( D => SIG_in(10), CK => clk, Q => n245
                           , QN => n_1058);
   MY_CLK_r_REG1121_S3 : DFF_X1 port map( D => SIG_in(9), CK => clk, Q => n244,
                           QN => n_1059);
   MY_CLK_r_REG1122_S3 : DFF_X1 port map( D => SIG_in(8), CK => clk, Q => n243,
                           QN => n_1060);
   MY_CLK_r_REG1135_S3 : DFF_X1 port map( D => SIG_in(7), CK => clk, Q => n242,
                           QN => n_1061);
   MY_CLK_r_REG1136_S3 : DFF_X1 port map( D => SIG_in(6), CK => clk, Q => n241,
                           QN => n_1062);
   MY_CLK_r_REG1138_S3 : DFF_X1 port map( D => SIG_in(5), CK => clk, Q => n240,
                           QN => n_1063);
   MY_CLK_r_REG1139_S3 : DFF_X1 port map( D => SIG_in(4), CK => clk, Q => 
                           n_1064, QN => n343);
   MY_CLK_r_REG1137_S3 : DFF_X1 port map( D => SIG_in(3), CK => clk, Q => n238,
                           QN => n337);
   MY_CLK_r_REG1152_S3 : DFF_X1 port map( D => SIG_in(2), CK => clk, Q => n237,
                           QN => n_1065);
   MY_CLK_r_REG1276_S1 : DFF_X1 port map( D => EXP_in(6), CK => clk, Q => 
                           n_1066, QN => n340);
   MY_CLK_r_REG1279_S1 : DFF_X1 port map( D => EXP_in(5), CK => clk, Q => 
                           n_1067, QN => n341);
   MY_CLK_r_REG1282_S1 : DFF_X1 port map( D => EXP_in(4), CK => clk, Q => 
                           n_1068, QN => n342);
   MY_CLK_r_REG1287_S3 : DFF_X1 port map( D => n231, CK => clk, Q => n230, QN 
                           => n344);
   MY_CLK_r_REG1296_S3 : DFF_X1 port map( D => n222, CK => clk, Q => n221, QN 
                           => n339);
   MY_CLK_r_REG1283_S2 : DFF_X1 port map( D => n342, CK => clk, Q => n220, QN 
                           => n_1069);
   MY_CLK_r_REG1284_S3 : DFF_X1 port map( D => n220, CK => clk, Q => n219, QN 
                           => n_1070);
   MY_CLK_r_REG1280_S2 : DFF_X1 port map( D => n341, CK => clk, Q => n218, QN 
                           => n_1071);
   MY_CLK_r_REG1281_S3 : DFF_X1 port map( D => n218, CK => clk, Q => n217, QN 
                           => n_1072);
   MY_CLK_r_REG1277_S2 : DFF_X1 port map( D => n340, CK => clk, Q => n216, QN 
                           => n_1073);
   MY_CLK_r_REG1278_S3 : DFF_X1 port map( D => n216, CK => clk, Q => n215, QN 
                           => n_1074);
   MY_CLK_r_REG1274_S2 : DFF_X1 port map( D => n338, CK => clk, Q => n214, QN 
                           => n_1075);
   MY_CLK_r_REG1275_S3 : DFF_X1 port map( D => n214, CK => clk, Q => n213, QN 
                           => n_1076);
   U56 : INV_X1 port map( A => SIG_in(27), ZN => n167);
   U14 : OR2_X1 port map( A1 => n344, A2 => n4, ZN => n162);
   U17 : BUF_X2 port map( A => SIG_in(27), Z => n345);
   MY_CLK_r_REG1273_S1 : DFF_X1 port map( D => EXP_in(7), CK => clk, Q => 
                           n_1077, QN => n338);
   MY_CLK_r_REG1295_S2 : DFF_X1 port map( D => n223, CK => clk, Q => n222, QN 
                           => n_1078);
   MY_CLK_r_REG1294_S1 : DFF_X1 port map( D => EXP_in(0), CK => clk, Q => n223,
                           QN => n_1079);
   MY_CLK_r_REG1293_S3 : DFF_X1 port map( D => n225, CK => clk, Q => n224, QN 
                           => n_1080);
   MY_CLK_r_REG1292_S2 : DFF_X1 port map( D => n226, CK => clk, Q => n225, QN 
                           => n_1081);
   MY_CLK_r_REG1291_S1 : DFF_X1 port map( D => EXP_in(1), CK => clk, Q => n226,
                           QN => n_1082);
   MY_CLK_r_REG1290_S3 : DFF_X1 port map( D => n228, CK => clk, Q => n227, QN 
                           => n_1083);
   MY_CLK_r_REG1289_S2 : DFF_X1 port map( D => n229, CK => clk, Q => n228, QN 
                           => n_1084);
   MY_CLK_r_REG1288_S1 : DFF_X1 port map( D => EXP_in(2), CK => clk, Q => n229,
                           QN => n_1085);
   MY_CLK_r_REG1286_S2 : DFF_X1 port map( D => n232, CK => clk, Q => n231, QN 
                           => n_1086);
   MY_CLK_r_REG1285_S1 : DFF_X1 port map( D => EXP_in(3), CK => clk, Q => n232,
                           QN => n_1087);
   U2 : CLKBUF_X2 port map( A => n345, Z => n52);

end SYN_FPnormalize;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage2_DW01_add_0 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic;  clk : in 
         std_logic);

end FPmul_stage2_DW01_add_0;

architecture SYN_rpl of FPmul_stage2_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port,
      carry_1_port, n2, n10, n11, n12, n13, n14 : std_logic;

begin
   
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => n2, S
                           => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U2 : XNOR2_X1 port map( A => B(0), B => A(0), ZN => SUM(0));
   U1 : OAI21_X1 port map( B1 => n12, B2 => n11, A => n10, ZN => carry_2_port);
   U3 : INV_X1 port map( A => carry_1_port, ZN => n12);
   U4 : OR2_X1 port map( A1 => B(0), A2 => A(0), ZN => carry_1_port);
   U5 : NOR2_X1 port map( A1 => B(1), A2 => A(1), ZN => n11);
   U6 : XNOR2_X1 port map( A => B(1), B => A(1), ZN => n13);
   U7 : NAND2_X1 port map( A1 => B(1), A2 => A(1), ZN => n10);
   U8 : XNOR2_X1 port map( A => carry_1_port, B => n13, ZN => SUM(1));
   U9 : XNOR2_X1 port map( A => n2, B => n14, ZN => SUM(7));
   U10 : XNOR2_X1 port map( A => A(7), B => B(7), ZN => n14);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity UnpackFP_1 is

   port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector 
         (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, isNaN,
         isINF, isZ, isDN : out std_logic);

end UnpackFP_1;

architecture SYN_UnpackFP of UnpackFP_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N13, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13_port, n14, 
      n29, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097 : 
      std_logic;

begin
   SIG <= ( n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, N13
      , FP(22), FP(21), FP(20), FP(19), FP(18), FP(17), FP(16), FP(15), FP(14),
      FP(13), FP(12), FP(11), FP(10), FP(9), FP(8), FP(7), FP(6), FP(5), FP(4),
      FP(3), FP(2), FP(1), FP(0) );
   EXP <= ( FP(30), FP(29), FP(28), FP(27), FP(26), FP(25), FP(24), FP(23) );
   SIGN <= FP(31);
   
   U19 : NAND3_X1 port map( A1 => n6, A2 => n7, A3 => n8, ZN => n2);
   U14 : NOR4_X1 port map( A1 => FP(18), A2 => FP(14), A3 => FP(16), A4 => 
                           FP(15), ZN => n6);
   U13 : NOR4_X1 port map( A1 => FP(11), A2 => FP(13), A3 => FP(12), A4 => 
                           FP(10), ZN => n7);
   U12 : NOR4_X1 port map( A1 => FP(8), A2 => FP(4), A3 => FP(6), A4 => FP(5), 
                           ZN => n9);
   U10 : NOR4_X1 port map( A1 => FP(21), A2 => FP(20), A3 => FP(17), A4 => 
                           FP(19), ZN => n11);
   U9 : NOR4_X1 port map( A1 => FP(22), A2 => FP(3), A3 => FP(2), A4 => FP(1), 
                           ZN => n12);
   U7 : NAND4_X1 port map( A1 => FP(26), A2 => FP(25), A3 => FP(24), A4 => 
                           FP(23), ZN => n4);
   U6 : NAND4_X1 port map( A1 => FP(30), A2 => FP(29), A3 => FP(28), A4 => 
                           FP(27), ZN => n5);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => isINF);
   U2 : NOR2_X1 port map( A1 => n2, A2 => N13, ZN => isZ);
   U3 : NOR2_X1 port map( A1 => n29, A2 => n3, ZN => isNaN);
   U17 : NOR4_X1 port map( A1 => FP(26), A2 => FP(25), A3 => FP(24), A4 => 
                           FP(23), ZN => n13_port);
   U16 : NOR4_X1 port map( A1 => FP(30), A2 => FP(29), A3 => FP(28), A4 => 
                           FP(27), ZN => n14);
   U5 : OR2_X1 port map( A1 => n4, A2 => n5, ZN => n3);
   U11 : INV_X1 port map( A => n2, ZN => n29);
   U18 : AND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n8)
                           ;
   U20 : NOR3_X1 port map( A1 => FP(0), A2 => FP(7), A3 => FP(9), ZN => n10);
   U8 : NAND2_X1 port map( A1 => n13_port, A2 => n14, ZN => N13);

end SYN_UnpackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity UnpackFP_0 is

   port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector 
         (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, isNaN,
         isINF, isZ, isDN : out std_logic);

end UnpackFP_0;

architecture SYN_UnpackFP of UnpackFP_0 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N13, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13_port, n14, 
      n15, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106 : 
      std_logic;

begin
   SIG <= ( n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, N13
      , FP(22), FP(21), FP(20), FP(19), FP(18), FP(17), FP(16), FP(15), FP(14),
      FP(13), FP(12), FP(11), FP(10), FP(9), FP(8), FP(7), FP(6), FP(5), FP(4),
      FP(3), FP(2), FP(1), FP(0) );
   EXP <= ( FP(30), FP(29), FP(28), FP(27), FP(26), FP(25), FP(24), FP(23) );
   SIGN <= FP(31);
   
   U19 : NAND3_X1 port map( A1 => n6, A2 => n7, A3 => n8, ZN => n2);
   U14 : NOR4_X1 port map( A1 => FP(18), A2 => FP(14), A3 => FP(16), A4 => 
                           FP(15), ZN => n6);
   U13 : NOR4_X1 port map( A1 => FP(11), A2 => FP(13), A3 => FP(12), A4 => 
                           FP(10), ZN => n7);
   U12 : NOR4_X1 port map( A1 => FP(8), A2 => FP(4), A3 => FP(6), A4 => FP(5), 
                           ZN => n9);
   U11 : NOR3_X1 port map( A1 => FP(0), A2 => FP(7), A3 => FP(9), ZN => n10);
   U10 : NOR4_X1 port map( A1 => FP(21), A2 => FP(20), A3 => FP(17), A4 => 
                           FP(19), ZN => n11);
   U9 : NOR4_X1 port map( A1 => FP(22), A2 => FP(3), A3 => FP(2), A4 => FP(1), 
                           ZN => n12);
   U7 : NAND4_X1 port map( A1 => FP(26), A2 => FP(25), A3 => FP(24), A4 => 
                           FP(23), ZN => n4);
   U6 : NAND4_X1 port map( A1 => FP(30), A2 => FP(29), A3 => FP(28), A4 => 
                           FP(27), ZN => n5);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => isINF);
   U3 : NOR2_X1 port map( A1 => n15, A2 => n3, ZN => isNaN);
   U8 : AND4_X1 port map( A1 => n9, A2 => n10, A3 => n11, A4 => n12, ZN => n8);
   U5 : OR2_X1 port map( A1 => n4, A2 => n5, ZN => n3);
   U2 : INV_X1 port map( A => n2, ZN => n15);
   U15 : NOR2_X1 port map( A1 => n2, A2 => N13, ZN => isZ);
   U18 : NAND2_X1 port map( A1 => n13_port, A2 => n14, ZN => N13);
   U16 : NOR4_X1 port map( A1 => FP(30), A2 => FP(29), A3 => FP(28), A4 => 
                           FP(27), ZN => n14);
   U17 : NOR4_X1 port map( A1 => FP(26), A2 => FP(25), A3 => FP(24), A4 => 
                           FP(23), ZN => n13_port);

end SYN_UnpackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage4 is

   port( EXP_neg : in std_logic;  EXP_out_round : in std_logic_vector (7 downto
         0);  EXP_pos, SIGN_out : in std_logic;  SIG_out_round : in 
         std_logic_vector (27 downto 0);  clk, isINF_tab, isNaN, isZ_tab : in 
         std_logic;  FP_Z : out std_logic_vector (31 downto 0));

end FPmul_stage4;

architecture SYN_struct of FPmul_stage4 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component PackFP
      port( SIGN : in std_logic;  EXP : in std_logic_vector (7 downto 0);  SIG 
            : in std_logic_vector (22 downto 0);  isNaN, isINF, isZ : in 
            std_logic;  FP : out std_logic_vector (31 downto 0);  clk : in 
            std_logic);
   end component;
   
   component FPnormalize_SIG_width28_1
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
            std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SIG_out_norm2_26_port, SIG_out_9_port, SIG_out_8_port, EXP_out_7_port
      , EXP_out_6_port, EXP_out_5_port, EXP_out_4_port, isINF, n12, n64, n151, 
      n152, n153, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n39,
      n46, n171, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n506, n389, n390, n391, n392, n393, n394, n395, n396, n398, 
      n400, n402, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
      n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, 
      n528, n529, n530, n531, n532, n533, n534, n535, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, 
      n_1132 : std_logic;

begin
   
   n151 <= '0';
   n152 <= '0';
   n153 <= '0';
   U18 : NAND3_X1 port map( A1 => n520, A2 => n514, A3 => n531, ZN => n10);
   U19 : NAND3_X1 port map( A1 => EXP_out_6_port, A2 => EXP_out_5_port, A3 => 
                           EXP_out_4_port, ZN => n15);
   U3 : NOR3_X1 port map( A1 => SIG_out_8_port, A2 => SIG_out_norm2_26_port, A3
                           => SIG_out_9_port, ZN => n12);
   U12 : NOR2_X1 port map( A1 => n515, A2 => n10, ZN => n4);
   U11 : NAND4_X1 port map( A1 => n510, A2 => n511, A3 => n509, A4 => n525, ZN 
                           => n6);
   U10 : NAND4_X1 port map( A1 => n526, A2 => n524, A3 => n507, A4 => n508, ZN 
                           => n7);
   U9 : NAND4_X1 port map( A1 => n530, A2 => n529, A3 => n512, A4 => n527, ZN 
                           => n8);
   U8 : NAND4_X1 port map( A1 => n532, A2 => n522, A3 => n528, A4 => n521, ZN 
                           => n9);
   U7 : NOR4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n5);
   U6 : NAND4_X1 port map( A1 => n513, A2 => n523, A3 => n4, A4 => n5, ZN => n3
                           );
   U16 : NOR2_X1 port map( A1 => n534, A2 => n15, ZN => n11);
   U4 : NOR2_X1 port map( A1 => EXP_out_7_port, A2 => n393, ZN => n14);
   U13 : INV_X1 port map( A => EXP_out_7_port, ZN => n171);
   U14 : AOI21_X1 port map( B1 => n11, B2 => n13, A => n14, ZN => n2);
   U17 : AOI21_X1 port map( B1 => n389, B2 => n2, A => n46, ZN => isINF);
   U15 : NOR4_X1 port map( A1 => n535, A2 => n39, A3 => n533, A4 => n171, ZN =>
                           n13);
   U5 : INV_X1 port map( A => n64, ZN => n39);
   U20 : OAI211_X1 port map( C1 => n395, C2 => n171, A => n391, B => n3, ZN => 
                           n46);
   MY_CLK_r_REG1065_S5 : DFF_X1 port map( D => n246, CK => clk, Q => n428, QN 
                           => n520);
   MY_CLK_r_REG1064_S5 : DFF_X1 port map( D => n245, CK => clk, Q => n427, QN 
                           => n521);
   MY_CLK_r_REG1063_S5 : DFF_X1 port map( D => n244, CK => clk, Q => n426, QN 
                           => n522);
   MY_CLK_r_REG1062_S5 : DFF_X1 port map( D => n243, CK => clk, Q => n425, QN 
                           => n523);
   MY_CLK_r_REG1061_S5 : DFF_X1 port map( D => n242, CK => clk, Q => n424, QN 
                           => n524);
   MY_CLK_r_REG1059_S5 : DFF_X1 port map( D => n241, CK => clk, Q => n423, QN 
                           => n525);
   MY_CLK_r_REG1058_S5 : DFF_X1 port map( D => n240, CK => clk, Q => n422, QN 
                           => n526);
   MY_CLK_r_REG1060_S5 : DFF_X1 port map( D => n239, CK => clk, Q => n421, QN 
                           => n527);
   MY_CLK_r_REG1071_S5 : DFF_X1 port map( D => n238, CK => clk, Q => n420, QN 
                           => n528);
   MY_CLK_r_REG1079_S5 : DFF_X1 port map( D => n237, CK => clk, Q => n419, QN 
                           => n529);
   MY_CLK_r_REG1055_S5 : DFF_X1 port map( D => n236, CK => clk, Q => n418, QN 
                           => n530);
   MY_CLK_r_REG1053_S5 : DFF_X1 port map( D => n235, CK => clk, Q => n417, QN 
                           => n531);
   MY_CLK_r_REG1051_S5 : DFF_X1 port map( D => n234, CK => clk, Q => n416, QN 
                           => n532);
   MY_CLK_r_REG1047_S5 : DFF_X1 port map( D => n233, CK => clk, Q => n415, QN 
                           => n507);
   MY_CLK_r_REG1076_S5 : DFF_X1 port map( D => n232, CK => clk, Q => n414, QN 
                           => n508);
   MY_CLK_r_REG1070_S5 : DFF_X1 port map( D => n231, CK => clk, Q => n413, QN 
                           => n509);
   MY_CLK_r_REG1078_S5 : DFF_X1 port map( D => n230, CK => clk, Q => n412, QN 
                           => n510);
   MY_CLK_r_REG1073_S5 : DFF_X1 port map( D => n229, CK => clk, Q => n411, QN 
                           => n511);
   MY_CLK_r_REG1075_S5 : DFF_X1 port map( D => n228, CK => clk, Q => n410, QN 
                           => n512);
   MY_CLK_r_REG1072_S5 : DFF_X1 port map( D => n227, CK => clk, Q => n409, QN 
                           => n513);
   MY_CLK_r_REG1074_S5 : DFF_X1 port map( D => n226, CK => clk, Q => n408, QN 
                           => n514);
   MY_CLK_r_REG1067_S5 : DFF_X1 port map( D => n225, CK => clk, Q => n407, QN 
                           => n534);
   MY_CLK_r_REG1077_S5 : DFF_X1 port map( D => n224, CK => clk, Q => n406, QN 
                           => n533);
   MY_CLK_r_REG1066_S5 : DFF_X1 port map( D => n223, CK => clk, Q => n405, QN 
                           => n535);
   MY_CLK_r_REG1270_S3 : DFF_X1 port map( D => n404, CK => clk, Q => n_1111, QN
                           => n516);
   MY_CLK_r_REG1265_S3 : DFF_X1 port map( D => n402, CK => clk, Q => n_1112, QN
                           => n517);
   MY_CLK_r_REG1026_S3 : DFF_X1 port map( D => n400, CK => clk, Q => n_1113, QN
                           => n518);
   MY_CLK_r_REG1036_S3 : DFF_X1 port map( D => n398, CK => clk, Q => n_1114, QN
                           => n519);
   MY_CLK_r_REG1045_S5 : DFF_X1 port map( D => n12, CK => clk, Q => n_1115, QN 
                           => n515);
   I1 : FPnormalize_SIG_width28_1 port map( SIG_in(27) => SIG_out_round(27), 
                           SIG_in(26) => SIG_out_round(26), SIG_in(25) => 
                           SIG_out_round(25), SIG_in(24) => SIG_out_round(24), 
                           SIG_in(23) => SIG_out_round(23), SIG_in(22) => 
                           SIG_out_round(22), SIG_in(21) => SIG_out_round(21), 
                           SIG_in(20) => SIG_out_round(20), SIG_in(19) => 
                           SIG_out_round(19), SIG_in(18) => SIG_out_round(18), 
                           SIG_in(17) => SIG_out_round(17), SIG_in(16) => 
                           SIG_out_round(16), SIG_in(15) => SIG_out_round(15), 
                           SIG_in(14) => SIG_out_round(14), SIG_in(13) => 
                           SIG_out_round(13), SIG_in(12) => SIG_out_round(12), 
                           SIG_in(11) => SIG_out_round(11), SIG_in(10) => 
                           SIG_out_round(10), SIG_in(9) => SIG_out_round(9), 
                           SIG_in(8) => SIG_out_round(8), SIG_in(7) => 
                           SIG_out_round(7), SIG_in(6) => SIG_out_round(6), 
                           SIG_in(5) => SIG_out_round(5), SIG_in(4) => 
                           SIG_out_round(4), SIG_in(3) => SIG_out_round(3), 
                           SIG_in(2) => n151, SIG_in(1) => n152, SIG_in(0) => 
                           n153, EXP_in(7) => EXP_out_round(7), EXP_in(6) => 
                           EXP_out_round(6), EXP_in(5) => EXP_out_round(5), 
                           EXP_in(4) => EXP_out_round(4), EXP_in(3) => 
                           EXP_out_round(3), EXP_in(2) => EXP_out_round(2), 
                           EXP_in(1) => EXP_out_round(1), EXP_in(0) => 
                           EXP_out_round(0), SIG_out(27) => n_1116, SIG_out(26)
                           => SIG_out_norm2_26_port, SIG_out(25) => n246, 
                           SIG_out(24) => n245, SIG_out(23) => n244, 
                           SIG_out(22) => n243, SIG_out(21) => n242, 
                           SIG_out(20) => n241, SIG_out(19) => n240, 
                           SIG_out(18) => n239, SIG_out(17) => n238, 
                           SIG_out(16) => n237, SIG_out(15) => n236, 
                           SIG_out(14) => n235, SIG_out(13) => n234, 
                           SIG_out(12) => SIG_out_9_port, SIG_out(11) => 
                           SIG_out_8_port, SIG_out(10) => n233, SIG_out(9) => 
                           n232, SIG_out(8) => n231, SIG_out(7) => n230, 
                           SIG_out(6) => n229, SIG_out(5) => n228, SIG_out(4) 
                           => n227, SIG_out(3) => n226, SIG_out(2) => n_1117, 
                           SIG_out(1) => n_1118, SIG_out(0) => n_1119, 
                           EXP_out(7) => EXP_out_7_port, EXP_out(6) => 
                           EXP_out_6_port, EXP_out(5) => EXP_out_5_port, 
                           EXP_out(4) => EXP_out_4_port, EXP_out(3) => n64, 
                           EXP_out(2) => n225, EXP_out(1) => n224, EXP_out(0) 
                           => n223, clk => clk);
   I3 : PackFP port map( SIGN => SIGN_out, EXP(7) => EXP_out_7_port, EXP(6) => 
                           EXP_out_6_port, EXP(5) => EXP_out_5_port, EXP(4) => 
                           EXP_out_4_port, EXP(3) => n64, EXP(2) => n407, 
                           EXP(1) => n406, EXP(0) => n405, SIG(22) => n428, 
                           SIG(21) => n427, SIG(20) => n426, SIG(19) => n425, 
                           SIG(18) => n424, SIG(17) => n423, SIG(16) => n422, 
                           SIG(15) => n421, SIG(14) => n420, SIG(13) => n419, 
                           SIG(12) => n418, SIG(11) => n417, SIG(10) => n416, 
                           SIG(9) => SIG_out_9_port, SIG(8) => SIG_out_8_port, 
                           SIG(7) => n415, SIG(6) => n414, SIG(5) => n413, 
                           SIG(4) => n412, SIG(3) => n411, SIG(2) => n410, 
                           SIG(1) => n409, SIG(0) => n408, isNaN => isNaN, 
                           isINF => isINF, isZ => n46, FP(31) => n506, FP(30) 
                           => FP_Z(30), FP(29) => FP_Z(29), FP(28) => FP_Z(28),
                           FP(27) => FP_Z(27), FP(26) => FP_Z(26), FP(25) => 
                           FP_Z(25), FP(24) => FP_Z(24), FP(23) => FP_Z(23), 
                           FP(22) => FP_Z(22), FP(21) => FP_Z(21), FP(20) => 
                           FP_Z(20), FP(19) => FP_Z(19), FP(18) => FP_Z(18), 
                           FP(17) => FP_Z(17), FP(16) => FP_Z(16), FP(15) => 
                           FP_Z(15), FP(14) => FP_Z(14), FP(13) => FP_Z(13), 
                           FP(12) => FP_Z(12), FP(11) => FP_Z(11), FP(10) => 
                           FP_Z(10), FP(9) => FP_Z(9), FP(8) => FP_Z(8), FP(7) 
                           => FP_Z(7), FP(6) => FP_Z(6), FP(5) => FP_Z(5), 
                           FP(4) => FP_Z(4), FP(3) => FP_Z(3), FP(2) => FP_Z(2)
                           , FP(1) => FP_Z(1), FP(0) => FP_Z(0), clk => clk);
   MY_CLK_r_REG1272_S5 : DFF_X1 port map( D => n396, CK => clk, Q => n395, QN 
                           => n_1120);
   MY_CLK_r_REG1271_S4 : DFF_X1 port map( D => n516, CK => clk, Q => n396, QN 
                           => n_1121);
   MY_CLK_r_REG1269_S2 : DFF_X1 port map( D => EXP_neg, CK => clk, Q => n404, 
                           QN => n_1122);
   MY_CLK_r_REG1267_S5 : DFF_X1 port map( D => n394, CK => clk, Q => n393, QN 
                           => n_1123);
   MY_CLK_r_REG1266_S4 : DFF_X1 port map( D => n517, CK => clk, Q => n394, QN 
                           => n_1124);
   MY_CLK_r_REG1264_S2 : DFF_X1 port map( D => EXP_pos, CK => clk, Q => n402, 
                           QN => n_1125);
   MY_CLK_r_REG1038_S5 : DFF_X1 port map( D => n392, CK => clk, Q => n391, QN 
                           => n_1126);
   MY_CLK_r_REG1037_S4 : DFF_X1 port map( D => n519, CK => clk, Q => n392, QN 
                           => n_1127);
   MY_CLK_r_REG1035_S2 : DFF_X1 port map( D => isZ_tab, CK => clk, Q => n398, 
                           QN => n_1128);
   MY_CLK_r_REG1028_S5 : DFF_X1 port map( D => n390, CK => clk, Q => n389, QN 
                           => n_1129);
   MY_CLK_r_REG1027_S4 : DFF_X1 port map( D => n518, CK => clk, Q => n390, QN 
                           => n_1130);
   MY_CLK_r_REG1025_S2 : DFF_X1 port map( D => isINF_tab, CK => clk, Q => n400,
                           QN => n_1131);
   MY_CLK_r_REG1020_S2 : DFF_X1 port map( D => n506, CK => clk, Q => FP_Z(31), 
                           QN => n_1132);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage3 is

   port( EXP_in : in std_logic_vector (7 downto 0);  EXP_neg_stage2, 
         EXP_pos_stage2, SIGN_out_stage2 : in std_logic;  SIG_in : in 
         std_logic_vector (27 downto 0);  clk, isINF_stage2, isNaN_stage2, 
         isZ_tab_stage2 : in std_logic;  EXP_neg : out std_logic;  
         EXP_out_round : out std_logic_vector (7 downto 0);  EXP_pos, SIGN_out 
         : out std_logic;  SIG_out_round : out std_logic_vector (27 downto 0); 
         isINF_tab, isNaN, isZ_tab : out std_logic);

end FPmul_stage3;

architecture SYN_struct of FPmul_stage3 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FPround_SIG_width28
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
            std_logic);
   end component;
   
   component FPnormalize_SIG_width28_0
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
            std_logic);
   end component;
   
   signal SIG_out_norm_27_port, SIG_out_norm_26_port, SIG_out_norm_25_port, 
      SIG_out_norm_24_port, SIG_out_norm_23_port, SIG_out_norm_22_port, 
      SIG_out_norm_21_port, SIG_out_norm_20_port, SIG_out_norm_19_port, 
      SIG_out_norm_18_port, SIG_out_norm_17_port, SIG_out_norm_16_port, 
      SIG_out_norm_15_port, SIG_out_norm_14_port, SIG_out_norm_13_port, 
      SIG_out_norm_12_port, SIG_out_norm_11_port, SIG_out_norm_10_port, 
      SIG_out_norm_9_port, SIG_out_norm_8_port, SIG_out_norm_7_port, 
      SIG_out_norm_6_port, SIG_out_norm_5_port, EXP_out_norm_7_port, 
      EXP_out_norm_6_port, EXP_out_norm_5_port, EXP_out_norm_4_port, 
      EXP_out_norm_3_port, EXP_out_norm_2_port, EXP_out_norm_1_port, 
      EXP_out_norm_0_port, n99, n100, n101, n102, n147, n149, n175, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149 : std_logic;

begin
   
   SIG_out_norm_27_port <= '0';
   n99 <= '0';
   n100 <= '0';
   n101 <= '0';
   n102 <= '0';
   I9 : FPnormalize_SIG_width28_0 port map( SIG_in(27) => SIG_in(27), 
                           SIG_in(26) => SIG_in(26), SIG_in(25) => SIG_in(25), 
                           SIG_in(24) => SIG_in(24), SIG_in(23) => SIG_in(23), 
                           SIG_in(22) => SIG_in(22), SIG_in(21) => SIG_in(21), 
                           SIG_in(20) => SIG_in(20), SIG_in(19) => SIG_in(19), 
                           SIG_in(18) => SIG_in(18), SIG_in(17) => SIG_in(17), 
                           SIG_in(16) => SIG_in(16), SIG_in(15) => SIG_in(15), 
                           SIG_in(14) => SIG_in(14), SIG_in(13) => SIG_in(13), 
                           SIG_in(12) => SIG_in(12), SIG_in(11) => SIG_in(11), 
                           SIG_in(10) => SIG_in(10), SIG_in(9) => SIG_in(9), 
                           SIG_in(8) => SIG_in(8), SIG_in(7) => SIG_in(7), 
                           SIG_in(6) => SIG_in(6), SIG_in(5) => SIG_in(5), 
                           SIG_in(4) => SIG_in(4), SIG_in(3) => SIG_in(3), 
                           SIG_in(2) => SIG_in(2), SIG_in(1) => n99, SIG_in(0) 
                           => n100, EXP_in(7) => EXP_in(7), EXP_in(6) => 
                           EXP_in(6), EXP_in(5) => EXP_in(5), EXP_in(4) => 
                           EXP_in(4), EXP_in(3) => EXP_in(3), EXP_in(2) => 
                           EXP_in(2), EXP_in(1) => EXP_in(1), EXP_in(0) => 
                           EXP_in(0), SIG_out(27) => n_1138, SIG_out(26) => 
                           SIG_out_norm_26_port, SIG_out(25) => 
                           SIG_out_norm_25_port, SIG_out(24) => 
                           SIG_out_norm_24_port, SIG_out(23) => 
                           SIG_out_norm_23_port, SIG_out(22) => 
                           SIG_out_norm_22_port, SIG_out(21) => 
                           SIG_out_norm_21_port, SIG_out(20) => 
                           SIG_out_norm_20_port, SIG_out(19) => 
                           SIG_out_norm_19_port, SIG_out(18) => 
                           SIG_out_norm_18_port, SIG_out(17) => 
                           SIG_out_norm_17_port, SIG_out(16) => 
                           SIG_out_norm_16_port, SIG_out(15) => 
                           SIG_out_norm_15_port, SIG_out(14) => 
                           SIG_out_norm_14_port, SIG_out(13) => 
                           SIG_out_norm_13_port, SIG_out(12) => 
                           SIG_out_norm_12_port, SIG_out(11) => 
                           SIG_out_norm_11_port, SIG_out(10) => 
                           SIG_out_norm_10_port, SIG_out(9) => 
                           SIG_out_norm_9_port, SIG_out(8) => 
                           SIG_out_norm_8_port, SIG_out(7) => 
                           SIG_out_norm_7_port, SIG_out(6) => 
                           SIG_out_norm_6_port, SIG_out(5) => 
                           SIG_out_norm_5_port, SIG_out(4) => n149, SIG_out(3) 
                           => n175, SIG_out(2) => n147, SIG_out(1) => n_1139, 
                           SIG_out(0) => n_1140, EXP_out(7) => 
                           EXP_out_norm_7_port, EXP_out(6) => 
                           EXP_out_norm_6_port, EXP_out(5) => 
                           EXP_out_norm_5_port, EXP_out(4) => 
                           EXP_out_norm_4_port, EXP_out(3) => 
                           EXP_out_norm_3_port, EXP_out(2) => 
                           EXP_out_norm_2_port, EXP_out(1) => 
                           EXP_out_norm_1_port, EXP_out(0) => 
                           EXP_out_norm_0_port, clk => clk);
   I11 : FPround_SIG_width28 port map( SIG_in(27) => SIG_out_norm_27_port, 
                           SIG_in(26) => SIG_out_norm_26_port, SIG_in(25) => 
                           SIG_out_norm_25_port, SIG_in(24) => 
                           SIG_out_norm_24_port, SIG_in(23) => 
                           SIG_out_norm_23_port, SIG_in(22) => 
                           SIG_out_norm_22_port, SIG_in(21) => 
                           SIG_out_norm_21_port, SIG_in(20) => 
                           SIG_out_norm_20_port, SIG_in(19) => 
                           SIG_out_norm_19_port, SIG_in(18) => 
                           SIG_out_norm_18_port, SIG_in(17) => 
                           SIG_out_norm_17_port, SIG_in(16) => 
                           SIG_out_norm_16_port, SIG_in(15) => 
                           SIG_out_norm_15_port, SIG_in(14) => 
                           SIG_out_norm_14_port, SIG_in(13) => 
                           SIG_out_norm_13_port, SIG_in(12) => 
                           SIG_out_norm_12_port, SIG_in(11) => 
                           SIG_out_norm_11_port, SIG_in(10) => 
                           SIG_out_norm_10_port, SIG_in(9) => 
                           SIG_out_norm_9_port, SIG_in(8) => 
                           SIG_out_norm_8_port, SIG_in(7) => 
                           SIG_out_norm_7_port, SIG_in(6) => 
                           SIG_out_norm_6_port, SIG_in(5) => 
                           SIG_out_norm_5_port, SIG_in(4) => n149, SIG_in(3) =>
                           n175, SIG_in(2) => n147, SIG_in(1) => n101, 
                           SIG_in(0) => n102, EXP_in(7) => EXP_out_norm_7_port,
                           EXP_in(6) => EXP_out_norm_6_port, EXP_in(5) => 
                           EXP_out_norm_5_port, EXP_in(4) => 
                           EXP_out_norm_4_port, EXP_in(3) => 
                           EXP_out_norm_3_port, EXP_in(2) => 
                           EXP_out_norm_2_port, EXP_in(1) => 
                           EXP_out_norm_1_port, EXP_in(0) => 
                           EXP_out_norm_0_port, SIG_out(27) => 
                           SIG_out_round(27), SIG_out(26) => SIG_out_round(26),
                           SIG_out(25) => SIG_out_round(25), SIG_out(24) => 
                           SIG_out_round(24), SIG_out(23) => SIG_out_round(23),
                           SIG_out(22) => SIG_out_round(22), SIG_out(21) => 
                           SIG_out_round(21), SIG_out(20) => SIG_out_round(20),
                           SIG_out(19) => SIG_out_round(19), SIG_out(18) => 
                           SIG_out_round(18), SIG_out(17) => SIG_out_round(17),
                           SIG_out(16) => SIG_out_round(16), SIG_out(15) => 
                           SIG_out_round(15), SIG_out(14) => SIG_out_round(14),
                           SIG_out(13) => SIG_out_round(13), SIG_out(12) => 
                           SIG_out_round(12), SIG_out(11) => SIG_out_round(11),
                           SIG_out(10) => SIG_out_round(10), SIG_out(9) => 
                           SIG_out_round(9), SIG_out(8) => SIG_out_round(8), 
                           SIG_out(7) => SIG_out_round(7), SIG_out(6) => 
                           SIG_out_round(6), SIG_out(5) => SIG_out_round(5), 
                           SIG_out(4) => SIG_out_round(4), SIG_out(3) => 
                           SIG_out_round(3), SIG_out(2) => n_1141, SIG_out(1) 
                           => n_1142, SIG_out(0) => n_1143, EXP_out(7) => 
                           EXP_out_round(7), EXP_out(6) => EXP_out_round(6), 
                           EXP_out(5) => EXP_out_round(5), EXP_out(4) => 
                           EXP_out_round(4), EXP_out(3) => EXP_out_round(3), 
                           EXP_out(2) => EXP_out_round(2), EXP_out(1) => 
                           EXP_out_round(1), EXP_out(0) => EXP_out_round(0), 
                           clk => clk);
   MY_CLK_r_REG1268_S1 : DFF_X1 port map( D => EXP_neg_stage2, CK => clk, Q => 
                           EXP_neg, QN => n_1144);
   MY_CLK_r_REG1263_S1 : DFF_X1 port map( D => EXP_pos_stage2, CK => clk, Q => 
                           EXP_pos, QN => n_1145);
   MY_CLK_r_REG1034_S1 : DFF_X1 port map( D => isZ_tab_stage2, CK => clk, Q => 
                           isZ_tab, QN => n_1146);
   MY_CLK_r_REG1029_S1 : DFF_X1 port map( D => isNaN_stage2, CK => clk, Q => 
                           isNaN, QN => n_1147);
   MY_CLK_r_REG1024_S1 : DFF_X1 port map( D => isINF_stage2, CK => clk, Q => 
                           isINF_tab, QN => n_1148);
   MY_CLK_r_REG1019_S1 : DFF_X1 port map( D => SIGN_out_stage2, CK => clk, Q =>
                           SIGN_out, QN => n_1149);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage2 is

   port( A_EXP : in std_logic_vector (7 downto 0);  A_SIG : in std_logic_vector
         (31 downto 0);  B_EXP : in std_logic_vector (7 downto 0);  B_SIG : in 
         std_logic_vector (31 downto 0);  SIGN_out_stage1, clk, isINF_stage1, 
         isNaN_stage1, isZ_tab_stage1 : in std_logic;  EXP_in : out 
         std_logic_vector (7 downto 0);  EXP_neg_stage2, EXP_pos_stage2, 
         SIGN_out_stage2 : out std_logic;  SIG_in : out std_logic_vector (27 
         downto 0);  isINF_stage2, isNaN_stage2, isZ_tab_stage2 : out std_logic
         );

end FPmul_stage2;

architecture SYN_struct of FPmul_stage2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X2
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component FPmul_stage2_DW01_add_0
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X4
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal mw_I4sum_7_port, n1, n19, n20, n21, n22, n23, n24, n25, 
      mult_143_n6630, mult_143_n6629, mult_143_n6628, mult_143_n6627, 
      mult_143_n6626, mult_143_n6625, mult_143_n6624, mult_143_n6621, 
      mult_143_n6620, mult_143_n6619, mult_143_n6611, mult_143_n6610, 
      mult_143_n6607, mult_143_n6605, mult_143_n6598, mult_143_n6597, 
      mult_143_n6592, mult_143_n6590, mult_143_n6589, mult_143_n6583, 
      mult_143_n6582, mult_143_n6581, mult_143_n6580, mult_143_n6578, 
      mult_143_n6577, mult_143_n6573, mult_143_n6572, mult_143_n6570, 
      mult_143_n6564, mult_143_n6563, mult_143_n6560, mult_143_n6559, 
      mult_143_n6555, mult_143_n6554, mult_143_n6551, mult_143_n6550, 
      mult_143_n6549, mult_143_n6543, mult_143_n6541, mult_143_n6536, 
      mult_143_n6535, mult_143_n6532, mult_143_n6526, mult_143_n6524, 
      mult_143_n6523, mult_143_n6518, mult_143_n6517, mult_143_n6516, 
      mult_143_n6513, mult_143_n6510, mult_143_n6501, mult_143_n6499, 
      mult_143_n6498, mult_143_n6496, mult_143_n6491, mult_143_n6490, 
      mult_143_n6479, mult_143_n6478, mult_143_n6473, mult_143_n6435, 
      mult_143_n6434, mult_143_n6432, mult_143_n6427, mult_143_n6421, 
      mult_143_n6417, mult_143_n6408, mult_143_n6407, mult_143_n6406, 
      mult_143_n6402, mult_143_n6401, mult_143_n6398, mult_143_n6397, 
      mult_143_n6388, mult_143_n6385, mult_143_n6382, mult_143_n6381, 
      mult_143_n6379, mult_143_n6374, mult_143_n6369, mult_143_n6368, 
      mult_143_n6367, mult_143_n6365, mult_143_n6362, mult_143_n6361, 
      mult_143_n6360, mult_143_n6348, mult_143_n6347, mult_143_n6346, 
      mult_143_n6322, mult_143_n6309, mult_143_n6308, mult_143_n6307, 
      mult_143_n6306, mult_143_n6305, mult_143_n6304, mult_143_n6303, 
      mult_143_n6302, mult_143_n6301, mult_143_n6300, mult_143_n6299, 
      mult_143_n6298, mult_143_n6297, mult_143_n6296, mult_143_n6295, 
      mult_143_n6294, mult_143_n6293, mult_143_n6292, mult_143_n6291, 
      mult_143_n6290, mult_143_n6289, mult_143_n6288, mult_143_n6287, 
      mult_143_n6286, mult_143_n6285, mult_143_n6284, mult_143_n6283, 
      mult_143_n6282, mult_143_n6279, mult_143_n6277, mult_143_n6276, 
      mult_143_n6275, mult_143_n6274, mult_143_n6273, mult_143_n6272, 
      mult_143_n6270, mult_143_n6269, mult_143_n6268, mult_143_n6267, 
      mult_143_n6266, mult_143_n6265, mult_143_n6264, mult_143_n6263, 
      mult_143_n6261, mult_143_n6260, mult_143_n6259, mult_143_n6258, 
      mult_143_n6257, mult_143_n6256, mult_143_n6255, mult_143_n6254, 
      mult_143_n6253, mult_143_n6252, mult_143_n6251, mult_143_n6250, 
      mult_143_n6249, mult_143_n6248, mult_143_n6247, mult_143_n6246, 
      mult_143_n6245, mult_143_n6244, mult_143_n6243, mult_143_n6242, 
      mult_143_n6241, mult_143_n6240, mult_143_n6239, mult_143_n6234, 
      mult_143_n6233, mult_143_n6232, mult_143_n6231, mult_143_n6230, 
      mult_143_n6229, mult_143_n6228, mult_143_n6226, mult_143_n6223, 
      mult_143_n6222, mult_143_n6219, mult_143_n6218, mult_143_n6217, 
      mult_143_n6216, mult_143_n6212, mult_143_n6210, mult_143_n6209, 
      mult_143_n6208, mult_143_n6207, mult_143_n6206, mult_143_n6205, 
      mult_143_n6204, mult_143_n6203, mult_143_n6201, mult_143_n6200, 
      mult_143_n6199, mult_143_n6198, mult_143_n6197, mult_143_n6196, 
      mult_143_n6195, mult_143_n6194, mult_143_n6193, mult_143_n6192, 
      mult_143_n6191, mult_143_n6190, mult_143_n6189, mult_143_n6186, 
      mult_143_n6184, mult_143_n6183, mult_143_n6182, mult_143_n6181, 
      mult_143_n6180, mult_143_n6179, mult_143_n6174, mult_143_n6173, 
      mult_143_n6172, mult_143_n6171, mult_143_n6170, mult_143_n6169, 
      mult_143_n6168, mult_143_n6167, mult_143_n6166, mult_143_n6165, 
      mult_143_n6162, mult_143_n6160, mult_143_n6159, mult_143_n6158, 
      mult_143_n6157, mult_143_n6156, mult_143_n6155, mult_143_n6154, 
      mult_143_n6149, mult_143_n6148, mult_143_n6147, mult_143_n6146, 
      mult_143_n6145, mult_143_n6144, mult_143_n6143, mult_143_n6142, 
      mult_143_n6141, mult_143_n6140, mult_143_n6139, mult_143_n6138, 
      mult_143_n6137, mult_143_n6136, mult_143_n6135, mult_143_n6134, 
      mult_143_n6133, mult_143_n6132, mult_143_n6131, mult_143_n6130, 
      mult_143_n6129, mult_143_n6128, mult_143_n6127, mult_143_n6126, 
      mult_143_n6125, mult_143_n6124, mult_143_n6123, mult_143_n6122, 
      mult_143_n6120, mult_143_n6119, mult_143_n6118, mult_143_n6115, 
      mult_143_n6114, mult_143_n6113, mult_143_n6112, mult_143_n6111, 
      mult_143_n6110, mult_143_n6109, mult_143_n6106, mult_143_n6105, 
      mult_143_n6104, mult_143_n6103, mult_143_n6102, mult_143_n6101, 
      mult_143_n6100, mult_143_n6099, mult_143_n6098, mult_143_n6097, 
      mult_143_n6096, mult_143_n6095, mult_143_n6093, mult_143_n6092, 
      mult_143_n6089, mult_143_n6088, mult_143_n6087, mult_143_n6086, 
      mult_143_n6085, mult_143_n6083, mult_143_n6082, mult_143_n6081, 
      mult_143_n6080, mult_143_n6079, mult_143_n6078, mult_143_n6076, 
      mult_143_n6075, mult_143_n6074, mult_143_n6073, mult_143_n6072, 
      mult_143_n6071, mult_143_n6070, mult_143_n6069, mult_143_n6068, 
      mult_143_n6067, mult_143_n6066, mult_143_n6065, mult_143_n6064, 
      mult_143_n6063, mult_143_n6062, mult_143_n6061, mult_143_n6059, 
      mult_143_n6058, mult_143_n6057, mult_143_n6056, mult_143_n6055, 
      mult_143_n6054, mult_143_n6053, mult_143_n6052, mult_143_n6051, 
      mult_143_n6050, mult_143_n6049, mult_143_n6048, mult_143_n6047, 
      mult_143_n6045, mult_143_n6043, mult_143_n6042, mult_143_n6041, 
      mult_143_n6040, mult_143_n6039, mult_143_n6038, mult_143_n6037, 
      mult_143_n6036, mult_143_n6035, mult_143_n6034, mult_143_n6033, 
      mult_143_n6031, mult_143_n6030, mult_143_n6029, mult_143_n6028, 
      mult_143_n6027, mult_143_n6026, mult_143_n6025, mult_143_n6024, 
      mult_143_n6023, mult_143_n6022, mult_143_n6020, mult_143_n6019, 
      mult_143_n6018, mult_143_n6017, mult_143_n6016, mult_143_n6015, 
      mult_143_n6014, mult_143_n6013, mult_143_n6012, mult_143_n6011, 
      mult_143_n6010, mult_143_n6009, mult_143_n6008, mult_143_n6005, 
      mult_143_n6004, mult_143_n6003, mult_143_n6002, mult_143_n6001, 
      mult_143_n6000, mult_143_n5999, mult_143_n5998, mult_143_n5997, 
      mult_143_n5995, mult_143_n5994, mult_143_n5992, mult_143_n5991, 
      mult_143_n5989, mult_143_n5988, mult_143_n5987, mult_143_n5986, 
      mult_143_n5985, mult_143_n5984, mult_143_n5982, mult_143_n5981, 
      mult_143_n5979, mult_143_n5978, mult_143_n5976, mult_143_n5975, 
      mult_143_n5974, mult_143_n5972, mult_143_n5971, mult_143_n5970, 
      mult_143_n5969, mult_143_n5967, mult_143_n5966, mult_143_n5965, 
      mult_143_n5964, mult_143_n5963, mult_143_n5962, mult_143_n5961, 
      mult_143_n5960, mult_143_n5959, mult_143_n5958, mult_143_n5956, 
      mult_143_n5955, mult_143_n5953, mult_143_n5952, mult_143_n5951, 
      mult_143_n5950, mult_143_n5949, mult_143_n5948, mult_143_n5946, 
      mult_143_n5945, mult_143_n5944, mult_143_n5943, mult_143_n5940, 
      mult_143_n5939, mult_143_n5938, mult_143_n5937, mult_143_n5936, 
      mult_143_n5935, mult_143_n5934, mult_143_n5933, mult_143_n5932, 
      mult_143_n5931, mult_143_n5930, mult_143_n5929, mult_143_n5928, 
      mult_143_n5927, mult_143_n5926, mult_143_n5925, mult_143_n5924, 
      mult_143_n5923, mult_143_n5922, mult_143_n5921, mult_143_n5920, 
      mult_143_n5919, mult_143_n5918, mult_143_n5917, mult_143_n5916, 
      mult_143_n5914, mult_143_n5913, mult_143_n5912, mult_143_n5910, 
      mult_143_n5907, mult_143_n5906, mult_143_n5905, mult_143_n5904, 
      mult_143_n5903, mult_143_n5901, mult_143_n5900, mult_143_n5899, 
      mult_143_n5898, mult_143_n5897, mult_143_n5896, mult_143_n5895, 
      mult_143_n5894, mult_143_n5893, mult_143_n5892, mult_143_n5889, 
      mult_143_n5888, mult_143_n5887, mult_143_n5886, mult_143_n5885, 
      mult_143_n5884, mult_143_n5883, mult_143_n5882, mult_143_n5881, 
      mult_143_n5880, mult_143_n5879, mult_143_n5878, mult_143_n5877, 
      mult_143_n5876, mult_143_n5875, mult_143_n5874, mult_143_n5873, 
      mult_143_n5872, mult_143_n5871, mult_143_n5870, mult_143_n5869, 
      mult_143_n5868, mult_143_n5867, mult_143_n5866, mult_143_n5865, 
      mult_143_n5864, mult_143_n5863, mult_143_n5862, mult_143_n5861, 
      mult_143_n5860, mult_143_n5859, mult_143_n5858, mult_143_n5857, 
      mult_143_n5855, mult_143_n5854, mult_143_n5853, mult_143_n5852, 
      mult_143_n5850, mult_143_n5849, mult_143_n5847, mult_143_n5846, 
      mult_143_n5845, mult_143_n5844, mult_143_n5842, mult_143_n5841, 
      mult_143_n5840, mult_143_n5837, mult_143_n5836, mult_143_n5834, 
      mult_143_n5833, mult_143_n5831, mult_143_n5830, mult_143_n5828, 
      mult_143_n5825, mult_143_n5824, mult_143_n5823, mult_143_n5822, 
      mult_143_n5821, mult_143_n5820, mult_143_n5819, mult_143_n5818, 
      mult_143_n5817, mult_143_n5816, mult_143_n5815, mult_143_n5814, 
      mult_143_n5813, mult_143_n5811, mult_143_n5810, mult_143_n5809, 
      mult_143_n5808, mult_143_n5807, mult_143_n5806, mult_143_n5805, 
      mult_143_n5804, mult_143_n5803, mult_143_n5802, mult_143_n5801, 
      mult_143_n5800, mult_143_n5799, mult_143_n5796, mult_143_n5794, 
      mult_143_n5793, mult_143_n5791, mult_143_n5789, mult_143_n5788, 
      mult_143_n5787, mult_143_n5786, mult_143_n5784, mult_143_n5783, 
      mult_143_n5782, mult_143_n5781, mult_143_n5780, mult_143_n5779, 
      mult_143_n5778, mult_143_n5777, mult_143_n5776, mult_143_n5775, 
      mult_143_n5772, mult_143_n5771, mult_143_n5770, mult_143_n5769, 
      mult_143_n5768, mult_143_n5765, mult_143_n5760, mult_143_n5758, 
      mult_143_n5755, mult_143_n5754, mult_143_n5751, mult_143_n5747, 
      mult_143_n5746, mult_143_n5743, mult_143_n5742, mult_143_n5741, 
      mult_143_n5740, mult_143_n5739, mult_143_n5738, mult_143_n5736, 
      mult_143_n5735, mult_143_n5733, mult_143_n5732, mult_143_n5731, 
      mult_143_n5730, mult_143_n5728, mult_143_n5725, mult_143_n5724, 
      mult_143_n5723, mult_143_n5722, mult_143_n5720, mult_143_n5719, 
      mult_143_n5718, mult_143_n5717, mult_143_n5716, mult_143_n5712, 
      mult_143_n5710, mult_143_n5709, mult_143_n5708, mult_143_n5707, 
      mult_143_n5706, mult_143_n5705, mult_143_n5704, mult_143_n5703, 
      mult_143_n5702, mult_143_n5701, mult_143_n5700, mult_143_n5699, 
      mult_143_n5698, mult_143_n5697, mult_143_n5696, mult_143_n5695, 
      mult_143_n5694, mult_143_n5693, mult_143_n5692, mult_143_n5691, 
      mult_143_n5690, mult_143_n5689, mult_143_n5688, mult_143_n5687, 
      mult_143_n5686, mult_143_n5685, mult_143_n5684, mult_143_n5683, 
      mult_143_n5682, mult_143_n5680, mult_143_n5679, mult_143_n5677, 
      mult_143_n5676, mult_143_n5673, mult_143_n5672, mult_143_n5671, 
      mult_143_n5670, mult_143_n5669, mult_143_n5668, mult_143_n5667, 
      mult_143_n5666, mult_143_n5665, mult_143_n5664, mult_143_n5663, 
      mult_143_n5662, mult_143_n5661, mult_143_n5660, mult_143_n5658, 
      mult_143_n5657, mult_143_n5656, mult_143_n5654, mult_143_n5653, 
      mult_143_n5652, mult_143_n5651, mult_143_n5650, mult_143_n5649, 
      mult_143_n5648, mult_143_n5647, mult_143_n5646, mult_143_n5643, 
      mult_143_n5641, mult_143_n5640, mult_143_n5639, mult_143_n5638, 
      mult_143_n5637, mult_143_n5636, mult_143_n5635, mult_143_n5634, 
      mult_143_n5633, mult_143_n5632, mult_143_n5631, mult_143_n5630, 
      mult_143_n5629, mult_143_n5628, mult_143_n5627, mult_143_n5626, 
      mult_143_n5625, mult_143_n5624, mult_143_n5623, mult_143_n5622, 
      mult_143_n5621, mult_143_n5620, mult_143_n5619, mult_143_n5618, 
      mult_143_n5617, mult_143_n5616, mult_143_n5615, mult_143_n5614, 
      mult_143_n5613, mult_143_n5612, mult_143_n5611, mult_143_n5610, 
      mult_143_n5609, mult_143_n5607, mult_143_n5606, mult_143_n5605, 
      mult_143_n5604, mult_143_n5601, mult_143_n5600, mult_143_n5598, 
      mult_143_n5597, mult_143_n5596, mult_143_n5595, mult_143_n5594, 
      mult_143_n5593, mult_143_n5592, mult_143_n5591, mult_143_n5590, 
      mult_143_n5589, mult_143_n5588, mult_143_n5587, mult_143_n5586, 
      mult_143_n5585, mult_143_n5583, mult_143_n5582, mult_143_n5581, 
      mult_143_n5580, mult_143_n5578, mult_143_n5576, mult_143_n5574, 
      mult_143_n5572, mult_143_n5571, mult_143_n5570, mult_143_n5569, 
      mult_143_n5568, mult_143_n5567, mult_143_n5566, mult_143_n5564, 
      mult_143_n5563, mult_143_n5562, mult_143_n5561, mult_143_n5559, 
      mult_143_n5558, mult_143_n5557, mult_143_n5556, mult_143_n5554, 
      mult_143_n5553, mult_143_n5552, mult_143_n5550, mult_143_n5547, 
      mult_143_n5545, mult_143_n5544, mult_143_n5543, mult_143_n5542, 
      mult_143_n5541, mult_143_n5540, mult_143_n5539, mult_143_n5534, 
      mult_143_n5533, mult_143_n5532, mult_143_n5531, mult_143_n5530, 
      mult_143_n5529, mult_143_n5528, mult_143_n5527, mult_143_n5526, 
      mult_143_n5525, mult_143_n5524, mult_143_n5523, mult_143_n5522, 
      mult_143_n5521, mult_143_n5517, mult_143_n5516, mult_143_n5515, 
      mult_143_n5514, mult_143_n5513, mult_143_n5512, mult_143_n5511, 
      mult_143_n5510, mult_143_n5509, mult_143_n5508, mult_143_n5507, 
      mult_143_n5505, mult_143_n5504, mult_143_n5503, mult_143_n5502, 
      mult_143_n5495, mult_143_n5494, mult_143_n5493, mult_143_n5492, 
      mult_143_n5491, mult_143_n5489, mult_143_n5488, mult_143_n5487, 
      mult_143_n5486, mult_143_n5485, mult_143_n5484, mult_143_n5483, 
      mult_143_n5481, mult_143_n5479, mult_143_n5478, mult_143_n5477, 
      mult_143_n5475, mult_143_n5474, mult_143_n5470, mult_143_n5469, 
      mult_143_n5468, mult_143_n5467, mult_143_n5466, mult_143_n5465, 
      mult_143_n5463, mult_143_n5462, mult_143_n5461, mult_143_n5456, 
      mult_143_n5450, mult_143_n5446, mult_143_n5445, mult_143_n5444, 
      mult_143_n5443, mult_143_n5441, mult_143_n5440, mult_143_n5439, 
      mult_143_n5437, mult_143_n5436, mult_143_n5435, mult_143_n5434, 
      mult_143_n5432, mult_143_n5431, mult_143_n5430, mult_143_n5426, 
      mult_143_n5425, mult_143_n5424, mult_143_n5422, mult_143_n5420, 
      mult_143_n5419, mult_143_n5418, mult_143_n5417, mult_143_n5416, 
      mult_143_n5415, mult_143_n5414, mult_143_n5413, mult_143_n5412, 
      mult_143_n5405, mult_143_n5404, mult_143_n5403, mult_143_n5402, 
      mult_143_n5401, mult_143_n5397, mult_143_n5396, mult_143_n5395, 
      mult_143_n5394, mult_143_n5393, mult_143_n5389, mult_143_n5387, 
      mult_143_n5385, mult_143_n5384, mult_143_n5382, mult_143_n5381, 
      mult_143_n5380, mult_143_n5379, mult_143_n5378, mult_143_n5377, 
      mult_143_n5376, mult_143_n5375, mult_143_n5374, mult_143_n5372, 
      mult_143_n5368, mult_143_n5367, mult_143_n5366, mult_143_n5365, 
      mult_143_n5363, mult_143_n5362, mult_143_n5361, mult_143_n5356, 
      mult_143_n5355, mult_143_n5354, mult_143_n5353, mult_143_n5352, 
      mult_143_n5351, mult_143_n5350, mult_143_n5347, mult_143_n5346, 
      mult_143_n5345, mult_143_n5344, mult_143_n5343, mult_143_n5342, 
      mult_143_n5341, mult_143_n5340, mult_143_n5338, mult_143_n5337, 
      mult_143_n5336, mult_143_n5335, mult_143_n5334, mult_143_n5333, 
      mult_143_n5332, mult_143_n5331, mult_143_n5330, mult_143_n5329, 
      mult_143_n5328, mult_143_n5327, mult_143_n5326, mult_143_n5325, 
      mult_143_n5324, mult_143_n5323, mult_143_n5322, mult_143_n5321, 
      mult_143_n5320, mult_143_n5318, mult_143_n5316, mult_143_n5315, 
      mult_143_n5313, mult_143_n5312, mult_143_n5311, mult_143_n5310, 
      mult_143_n5309, mult_143_n5307, mult_143_n5306, mult_143_n5305, 
      mult_143_n5304, mult_143_n5303, mult_143_n5300, mult_143_n5299, 
      mult_143_n5298, mult_143_n5297, mult_143_n5296, mult_143_n5294, 
      mult_143_n5293, mult_143_n5291, mult_143_n5290, mult_143_n5289, 
      mult_143_n5288, mult_143_n5285, mult_143_n5284, mult_143_n5280, 
      mult_143_n5279, mult_143_n5278, mult_143_n5276, mult_143_n5275, 
      mult_143_n5274, mult_143_n5273, mult_143_n5272, mult_143_n5271, 
      mult_143_n5270, mult_143_n5269, mult_143_n5268, mult_143_n5267, 
      mult_143_n5266, mult_143_n5265, mult_143_n5264, mult_143_n5263, 
      mult_143_n5262, mult_143_n5261, mult_143_n5260, mult_143_n5259, 
      mult_143_n5258, mult_143_n5257, mult_143_n5256, mult_143_n5255, 
      mult_143_n5254, mult_143_n5253, mult_143_n5252, mult_143_n5251, 
      mult_143_n5250, mult_143_n5243, mult_143_n5242, mult_143_n5240, 
      mult_143_n5239, mult_143_n5236, mult_143_n5235, mult_143_n5232, 
      mult_143_n5231, mult_143_n5230, mult_143_n5228, mult_143_n5221, 
      mult_143_n5219, mult_143_n5216, mult_143_n5215, mult_143_n5209, 
      mult_143_n5208, mult_143_n5207, mult_143_n5206, mult_143_n5205, 
      mult_143_n5204, mult_143_n5203, mult_143_n5201, mult_143_n5200, 
      mult_143_n5199, mult_143_n5197, mult_143_n5196, mult_143_n5195, 
      mult_143_n5194, mult_143_n5193, mult_143_n5192, mult_143_n5191, 
      mult_143_n5190, mult_143_n5189, mult_143_n5188, mult_143_n5187, 
      mult_143_n5186, mult_143_n5185, mult_143_n5184, mult_143_n5182, 
      mult_143_n5181, mult_143_n5180, mult_143_n5179, mult_143_n5178, 
      mult_143_n5177, mult_143_n5176, mult_143_n5175, mult_143_n5174, 
      mult_143_n5170, mult_143_n5169, mult_143_n5168, mult_143_n5166, 
      mult_143_n5165, mult_143_n5164, mult_143_n5163, mult_143_n5162, 
      mult_143_n5161, mult_143_n5160, mult_143_n5159, mult_143_n5158, 
      mult_143_n5153, mult_143_n5152, mult_143_n5145, mult_143_n5144, 
      mult_143_n5143, mult_143_n5142, mult_143_n5138, mult_143_n5137, 
      mult_143_n5136, mult_143_n5135, mult_143_n5134, mult_143_n5133, 
      mult_143_n5132, mult_143_n5131, mult_143_n5130, mult_143_n5129, 
      mult_143_n5128, mult_143_n5127, mult_143_n5126, mult_143_n5125, 
      mult_143_n5124, mult_143_n5123, mult_143_n5122, mult_143_n5121, 
      mult_143_n5120, mult_143_n5119, mult_143_n5118, mult_143_n5117, 
      mult_143_n5111, mult_143_n5095, mult_143_n5094, mult_143_n5092, 
      mult_143_n5090, mult_143_n5089, mult_143_n5087, mult_143_n5086, 
      mult_143_n5085, mult_143_n5084, mult_143_n5083, mult_143_n5080, 
      mult_143_n5075, mult_143_n5074, mult_143_n5071, mult_143_n5070, 
      mult_143_n5069, mult_143_n5068, mult_143_n5067, mult_143_n5065, 
      mult_143_n5059, mult_143_n5058, mult_143_n5057, mult_143_n5054, 
      mult_143_n5052, mult_143_n5050, mult_143_n5048, mult_143_n5047, 
      mult_143_n5046, mult_143_n5041, mult_143_n5040, mult_143_n5035, 
      mult_143_n5033, mult_143_n5028, mult_143_n5027, mult_143_n5025, 
      mult_143_n5023, mult_143_n5020, mult_143_n5019, mult_143_n5018, 
      mult_143_n5017, mult_143_n5016, mult_143_n5015, mult_143_n5012, 
      mult_143_n5009, mult_143_n5008, mult_143_n5007, mult_143_n5004, 
      mult_143_n5002, mult_143_n5001, mult_143_n4995, mult_143_n4994, 
      mult_143_n4991, mult_143_n4989, mult_143_n4988, mult_143_n4987, 
      mult_143_n4985, mult_143_n4984, mult_143_n4981, mult_143_n4980, 
      mult_143_n4973, mult_143_n4972, mult_143_n4971, mult_143_n4970, 
      mult_143_n4966, mult_143_n4965, mult_143_n4963, mult_143_n4962, 
      mult_143_n4961, mult_143_n4960, mult_143_n4959, mult_143_n4957, 
      mult_143_n4956, mult_143_n4954, mult_143_n4953, mult_143_n4949, 
      mult_143_n4948, mult_143_n4947, mult_143_n4946, mult_143_n4945, 
      mult_143_n4944, mult_143_n4943, mult_143_n4942, mult_143_n4941, 
      mult_143_n4939, mult_143_n4937, mult_143_n4936, mult_143_n4935, 
      mult_143_n4934, mult_143_n4933, mult_143_n4932, mult_143_n4931, 
      mult_143_n4928, mult_143_n4927, mult_143_n4926, mult_143_n4925, 
      mult_143_n4924, mult_143_n4923, mult_143_n4922, mult_143_n4920, 
      mult_143_n4919, mult_143_n4915, mult_143_n4914, mult_143_n4913, 
      mult_143_n4910, mult_143_n4909, mult_143_n4908, mult_143_n4905, 
      mult_143_n4903, mult_143_n4902, mult_143_n4901, mult_143_n4900, 
      mult_143_n4897, mult_143_n4896, mult_143_n4895, mult_143_n4894, 
      mult_143_n4893, mult_143_n4892, mult_143_n4891, mult_143_n4890, 
      mult_143_n4889, mult_143_n4888, mult_143_n4887, mult_143_n4886, 
      mult_143_n4883, mult_143_n4881, mult_143_n4880, mult_143_n4879, 
      mult_143_n4878, mult_143_n4877, mult_143_n4876, mult_143_n4875, 
      mult_143_n4874, mult_143_n4870, mult_143_n4869, mult_143_n4864, 
      mult_143_n4863, mult_143_n4862, mult_143_n4861, mult_143_n4860, 
      mult_143_n4859, mult_143_n4858, mult_143_n4857, mult_143_n4856, 
      mult_143_n4853, mult_143_n4852, mult_143_n4851, mult_143_n4850, 
      mult_143_n4849, mult_143_n4848, mult_143_n4846, mult_143_n4845, 
      mult_143_n4844, mult_143_n4843, mult_143_n4842, mult_143_n4841, 
      mult_143_n4840, mult_143_n4839, mult_143_n4838, mult_143_n4837, 
      mult_143_n4832, mult_143_n4831, mult_143_n4830, mult_143_n4829, 
      mult_143_n4828, mult_143_n4827, mult_143_n4826, mult_143_n4825, 
      mult_143_n4824, mult_143_n4823, mult_143_n4822, mult_143_n4821, 
      mult_143_n4820, mult_143_n4819, mult_143_n4818, mult_143_n4815, 
      mult_143_n4813, mult_143_n4812, mult_143_n4811, mult_143_n4810, 
      mult_143_n4809, mult_143_n4808, mult_143_n4807, mult_143_n4806, 
      mult_143_n4805, mult_143_n4804, mult_143_n4803, mult_143_n4802, 
      mult_143_n4801, mult_143_n4800, mult_143_n4799, mult_143_n4798, 
      mult_143_n4797, mult_143_n4796, mult_143_n4795, mult_143_n4794, 
      mult_143_n4793, mult_143_n4792, mult_143_n4791, mult_143_n4790, 
      mult_143_n4789, mult_143_n4788, mult_143_n4787, mult_143_n4786, 
      mult_143_n4785, mult_143_n4784, mult_143_n4783, mult_143_n4782, 
      mult_143_n4781, mult_143_n4780, mult_143_n4779, mult_143_n4778, 
      mult_143_n4777, mult_143_n4776, mult_143_n4775, mult_143_n4774, 
      mult_143_n4773, mult_143_n4771, mult_143_n4768, mult_143_n4767, 
      mult_143_n4766, mult_143_n4762, mult_143_n4761, mult_143_n4760, 
      mult_143_n4759, mult_143_n4758, mult_143_n4757, mult_143_n4756, 
      mult_143_n4755, mult_143_n4555, mult_143_n4510, mult_143_n4504, 
      mult_143_n4502, mult_143_n4493, mult_143_n4490, mult_143_n4475, 
      mult_143_n4468, mult_143_n4467, mult_143_n4407, mult_143_n4401, 
      mult_143_n4366, mult_143_n4363, mult_143_n4361, mult_143_n4359, 
      mult_143_n4357, mult_143_n4355, mult_143_n4351, mult_143_n4348, 
      mult_143_n4344, mult_143_n4340, mult_143_n4339, mult_143_n4327, 
      mult_143_n4325, mult_143_n4319, mult_143_n4317, mult_143_n4309, 
      mult_143_n4307, mult_143_n4301, mult_143_n4275, mult_143_n4273, 
      mult_143_n4217, mult_143_n4215, mult_143_n4208, mult_143_n4206, 
      mult_143_n4201, mult_143_n4199, mult_143_n4156, mult_143_n4154, 
      mult_143_n3455, mult_143_n3448, mult_143_n3443, mult_143_n1904, 
      mult_143_n777, mult_143_n96, mult_143_n335, mult_143_n344, mult_143_n276,
      mult_143_n2755, mult_143_n304, mult_143_n904, mult_143_n922, 
      mult_143_n364, mult_143_n373, mult_143_n2200, mult_143_n3245, 
      mult_143_n3239, mult_143_n3228, mult_143_n3154, mult_143_n3137, 
      mult_143_n3096, mult_143_n3094, mult_143_n3083, mult_143_n3075, 
      mult_143_n3073, mult_143_n3055, mult_143_n3010, mult_143_n3007, 
      mult_143_n2981, mult_143_n2919, mult_143_n2868, mult_143_n2800, 
      mult_143_n2798, mult_143_n2772, mult_143_n2759, mult_143_n2743, 
      mult_143_n2702, mult_143_n2458, mult_143_n2401, mult_143_n2334, 
      mult_143_n2267, mult_143_n2133, mult_143_n2066, mult_143_n2001, 
      mult_143_n1942, mult_143_n1912, mult_143_n1911, mult_143_n1910, 
      mult_143_n1909, mult_143_n1908, mult_143_n1907, mult_143_n1906, 
      mult_143_n1905, mult_143_n1902, mult_143_n1901, mult_143_n1900, 
      mult_143_n1898, mult_143_n1897, mult_143_n1896, mult_143_n1895, 
      mult_143_n1894, mult_143_n1893, mult_143_n1892, mult_143_n1891, 
      mult_143_n1863, mult_143_n1853, mult_143_n1818, mult_143_n1816, 
      mult_143_n1815, mult_143_n1754, mult_143_n1753, mult_143_n1724, 
      mult_143_n1719, mult_143_n1690, mult_143_n1610, mult_143_n1582, 
      mult_143_n1553, mult_143_n1537, mult_143_n1536, mult_143_n1532, 
      mult_143_n1530, mult_143_n1528, mult_143_n1523, mult_143_n1521, 
      mult_143_n1127, mult_143_n1123, mult_143_n1116, mult_143_n1101, 
      mult_143_n1070, mult_143_n1059, mult_143_n1039, mult_143_n1027, 
      mult_143_n1017, mult_143_n1005, mult_143_n994, mult_143_n977, 
      mult_143_n938, mult_143_n917, mult_143_n901, mult_143_n897, mult_143_n886
      , mult_143_n867, mult_143_n813, mult_143_n812, mult_143_n811, 
      mult_143_n809, mult_143_n795, mult_143_n759, mult_143_n744, mult_143_n724
      , mult_143_n706, mult_143_n686, mult_143_n671, mult_143_n655, 
      mult_143_n654, mult_143_n652, mult_143_n650, mult_143_n610, mult_143_n581
      , mult_143_n522, mult_143_n430, mult_143_n427, mult_143_n426, 
      mult_143_n412, mult_143_n405, mult_143_n393, mult_143_n392, mult_143_n218
      , mult_143_n84, mult_143_n76, mult_143_n74, mult_143_n72, mult_143_n48, 
      mult_143_n36, mult_143_n2, n378, n380, n381, n382, n385, n386, n387, n388
      , n391, n392, n394, n395, n396, n397, n398, n400, n403, n404, n407, n408,
      n413, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n431, n433, n434, n435, n436, n438, n440, n441, n442, n445, n446, 
      n453, n456, n457, n460, n461, n463, n464, n465, n471, n473, n478, n479, 
      n480, n482, n484, n485, n486, n487, n490, n493, n494, n496, n500, n501, 
      n505, n506, n507, n508, n511, n512, n513, n514, n515, n516, n518, n519, 
      n523, n525, n527, n528, n532, n533, n536, n537, n538, n539, n542, n544, 
      n545, n546, n547, n548, n549, n552, n553, n555, n557, n558, n560, n562, 
      n563, n564, n565, n566, n567, n568, n569, n571, n572, n573, n581, n582, 
      n583, n584, n585, n587, n595, n599, n601, n603, n604, n605, n606, n607, 
      n608, n611, n616, n617, n618, n620, n624, n629, n630, n631, n632, n633, 
      n634, n636, n637, n638, n639, n641, n642, n643, n646, n648, n649, n650, 
      n651, n654, n657, n660, n666, n667, n671, n680, n686, n688, n693, n698, 
      n699, n702, n711, n712, n714, n715, n716, n717, n718, n720, n721, n724, 
      n726, n727, n728, n730, n734, n740, n743, n744, n745, n747, n748, n755, 
      n765, n772, n774, n778, n787, n799, n804, n808, n809, n811, n812, n813, 
      n814, n816, n817, n818, n819, n820, n821, n824, n825, n826, n847, n851, 
      n852, n860, n865, n868, n874, n878, n882, n886, n891, n895, n909, n910, 
      n942, n943, n944, n945, n946, n948, n949, n951, n953, n954, n955, n956, 
      n957, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, 
      n972, n974, n975, n976, n977, n978, n979, n980, n981, n982, n984, n986, 
      n990, n991, n992, n993, n994, n996, n997, n1003, n1005, n1008, n1010, 
      n1011, n1013, n1018, n1019, n1023, n1024, n1026, n1027, n1030, n1031, 
      n1032, n1034, n1035, n1037, n1038, n1039, n1040, n1042, n1045, n1046, 
      n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1055, n1056, n1057, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1075, n1077, n1078, n1079, n1083, n1085, n1469, 
      n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
      n1480, n1481, n1482, n1483, n1484, n1486, n1488, n1489, n1490, n1491, 
      n1493, n1494, n1498, n1499, n1500, n1501, n1502, n1503, n1505, n1507, 
      n1508, n1514, n1515, n1516, n1517, n1520, n1521, n1522, n1523, n1524, 
      n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1541, n1542, n1543, n1544, n1545, n1547, 
      n1548, n1549, n1550, n1551, n1552, n1555, n1556, n1557, n1558, n1559, 
      n1560, n1561, n1562, n1563, n1564, n1565, n1567, n1568, n1570, n1571, 
      n1572, n1573, n1574, n1575, n1577, n1578, n1579, n1582, n1584, n1587, 
      n1588, n1589, n1590, n1594, n1596, n1597, n1600, n1601, n1604, n1606, 
      n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
      n1617, n1618, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
      n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, 
      n1638, n1639, n1640, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
      n1650, n1651, n1657, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1683, n1684, n1685, n1686, 
      n1687, n1688, n1689, n1691, n1693, n1695, n1697, n1698, n1699, n1700, 
      n1701, n1702, n1703, n1705, n1706, n1707, n1708, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1718, n1719, n1720, n1721, n1722, n1723, n1724, 
      n1725, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, 
      n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
      n1756, n1757, n1758, n1759, n1765, n1782, n1787, n1828, n1832, n1836, 
      n1839, n1840, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, 
      n2606, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2617, 
      n2618, n2619, n2620, n2621, n2622, n2624, n2627, n2630, n2631, n2632, 
      n2633, n2634, n2636, n2637, n2638, n2664, n2665, n2666, n2667, n2668, 
      n2669, n2670, n2672, n2675, n2679, n2685, n2686, n2688, n2689, n2690, 
      n2691, n2692, n2694, n2695, n2696, n2703, n2704, n2705, n2706, n2707, 
      n2709, n2710, n2711, n2713, n2714, n2715, n2716, n2717, n2718, n2719, 
      n2720, n2721, n2722, n2723, n2725, n2726, n2727, n2728, n2730, n2731, 
      n2732, n2733, n2736, n2737, n2739, n2746, n2747, n2749, n2750, n2751, 
      n2755, n2756, n2757, n2759, n2761, n2762, n2764, n2765, n2766, n2767, 
      n2768, n2769, n2770, n2778, n2780, n2782, n2784, n2786, n2791, n2792, 
      n2793, n2794, n2796, n2799, n2803, n2804, n2805, n2806, n2811, n2812, 
      n2814, n2817, n2823, n2824, n2825, n2829, n2830, n2831, n2835, n2837, 
      n2840, n2841, n2844, n2846, n2847, n2848, n2850, n2851, n2852, n2855, 
      n2859, n2861, n2864, n2865, n2869, n2874, n2875, n2877, n2881, n2884, 
      n2885, n2888, n2890, n2891, n2893, n2895, n2898, n2901, n2905, n2906, 
      n2908, n2909, n2910, n2911, n2913, n2918, n2920, n2922, n2923, n2924, 
      n2927, n2934, n2936, n2937, n2938, n2945, n2947, n2948, n2951, n2952, 
      n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2962, n2963, 
      n2964, n2966, n2967, n2970, n2971, n2972, n2973, n2974, n2975, n2976, 
      n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, 
      n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, 
      n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, 
      n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, 
      n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, 
      n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3036, n3037, 
      n3038, n3039, n3040, n3041, n3042, n3044, n3045, n3046, n3047, n3048, 
      n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, 
      n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, 
      n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, 
      n3079, n3080, n3082, n3083, n3084, n3085, n3086, n3087, n3090, n3091, 
      n3093, n3095, n3097, n3099, n3100, n3101, n3104, n3105, n3106, n3107, 
      n3108, n3110, n3112, n3115, n3116, n3117, n3118, n3120, n3121, n3122, 
      n3123, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, 
      n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, 
      n3508, n3509, n3510, n3511, n3512, n3513, n3515, n3516, n3517, n3518, 
      n3519, n3520, n3521, n3523, n3524, n3525, n3526, n3527, n3528, n3529, 
      n3530, n3531, n3532, n3533, n3535, n3536, n3537, n3538, n3539, n3540, 
      n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3551, n3552, 
      n3553, n3554, n3555, n3556, n3558, n3559, n3560, n3561, n3562, n3563, 
      n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, 
      n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, 
      n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, 
      n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, 
      n3605, n3606, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, 
      n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, 
      n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, 
      n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, 
      n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, 
      n3656, n3657, n3658, n3659, n3660, n3662, n3663, n3664, n3665, n3666, 
      n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, 
      n3677, n3678, n3680, n3681, n3682, n3683, n3685, n3686, n3687, n3688, 
      n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, 
      n3699, n3700, n3701, n3702, n3703, n3705, n3706, n3707, n3708, n3709, 
      n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, 
      n3721, n3722, n3723, n3724, n3725, n3726, n3728, n3729, n3730, n3731, 
      n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
      n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, 
      n3752, n3754, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, 
      n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, 
      n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, 
      n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, 
      n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, 
      n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, 
      n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, 
      n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n4567, n4568, 
      n4569, n4570, n4571, n4573, n4574, n4575, n4576, n4577, n4578, n4579, 
      n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, 
      n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, 
      n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, 
      n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, 
      n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, 
      n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, 
      n4640, n4641, n4642, n4644, n4645, n4646, n4647, n4648, n4649, n4650, 
      n4651, n4652, n4653, n4655, n4656, n4657, n4658, n4661, n4662, n4663, 
      n4664, n4665, n4667, n4669, n4670, n4671, n4672, n4673, n4674, n4675, 
      n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4685, n4686, 
      n4688, n4689, n4690, n4692, n4693, n4694, n4695, n4697, n4699, n4700, 
      n4701, n4702, n4703, n4704, n4709, n4710, n4713, n4714, n4716, n4717, 
      n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, 
      n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, 
      n4738, n4739, n4742, n4743, n4744, n4746, n4747, n4748, n4749, n4750, 
      n4751, n4752, n4753, n4754, n4755, n4756, n4758, n4759, n4760, n4761, 
      n4762, n4763, n4764, n4765, n4766, n4768, n4769, n4770, n4771, n4772, 
      n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, 
      n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4826, n4827, 
      n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, 
      n4838, n4839, n4841, n4842, n4843, n4844, n4845, n4847, n4848, n4849, 
      n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, 
      n4860, n4861, n4862, n4863, n4864, n4866, n4867, n4868, n4869, n4870, 
      n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, 
      n4882, n4883, n4885, n4886, n4887, n4888, n4889, n4890, n4892, n4894, 
      n4895, n4896, n4901, n4903, n4904, n4905, n4906, n4907, n4908, n4909, 
      n4910, n4912, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, 
      n4928, n4929, n4930, n4932, n4933, n4935, n4936, n4937, n4938, n4939, 
      n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4949, n4950, 
      n4951, n4952, n4955, n4956, n4963, n4964, n4965, n4966, n4967, n4968, 
      n4969, n4970, n4971, n4972, n4973, n4979, n4980, n4981, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, 
      n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, 
      n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, 
      n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, 
      n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, 
      n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415 : std_logic;

begin
   SIGN_out_stage2 <= SIGN_out_stage1;
   isINF_stage2 <= isINF_stage1;
   isNaN_stage2 <= isNaN_stage1;
   isZ_tab_stage2 <= isZ_tab_stage1;
   
   n1 <= '1';
   U42 : NAND3_X1 port map( A1 => B_EXP(5), A2 => B_EXP(0), A3 => B_EXP(1), ZN 
                           => n23);
   U43 : NAND3_X1 port map( A1 => A_EXP(5), A2 => A_EXP(0), A3 => A_EXP(1), ZN 
                           => n21);
   U40 : NAND4_X1 port map( A1 => A_EXP(2), A2 => A_EXP(3), A3 => A_EXP(6), A4 
                           => A_EXP(4), ZN => n20);
   U39 : NAND4_X1 port map( A1 => B_EXP(2), A2 => B_EXP(3), A3 => B_EXP(6), A4 
                           => B_EXP(4), ZN => n22);
   U38 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => n22, B2 => n23, ZN => 
                           n19);
   U37 : NOR3_X1 port map( A1 => B_EXP(7), A2 => A_EXP(7), A3 => n19, ZN => 
                           EXP_neg_stage2);
   U36 : NOR2_X1 port map( A1 => n24, A2 => n25, ZN => EXP_pos_stage2);
   mult_143_U3936 : XNOR2_X1 port map( A => n1765, B => A_SIG(10), ZN => 
                           mult_143_n6243);
   mult_143_U4011 : NOR2_X1 port map( A1 => n651, A2 => mult_143_n6301, ZN => 
                           mult_143_n76);
   mult_143_U3994 : XNOR2_X1 port map( A => n649, B => A_SIG(13), ZN => 
                           mult_143_n6284);
   mult_143_U2720 : AOI222_X1 port map( A1 => mult_143_n1853, A2 => 
                           mult_143_n5084, B1 => mult_143_n1853, B2 => n688, C1
                           => mult_143_n5084, C2 => n688, ZN => mult_143_n654);
   mult_143_U2718 : XNOR2_X1 port map( A => mult_143_n1853, B => mult_143_n5083
                           , ZN => mult_143_n655);
   mult_143_U2719 : AOI22_X1 port map( A1 => mult_143_n1815, A2 => n680, B1 => 
                           mult_143_n5084, B2 => n688, ZN => mult_143_n5083);
   mult_143_U2721 : AOI21_X1 port map( B1 => n1782, B2 => n1828, A => 
                           mult_143_n5085, ZN => mult_143_n5084);
   mult_143_U2722 : AOI21_X1 port map( B1 => A_SIG(8), B2 => mult_143_n1818, A 
                           => mult_143_n1816, ZN => mult_143_n5085);
   mult_143_U3734 : AOI222_X1 port map( A1 => mult_143_n4317, A2 => B_SIG(11), 
                           B1 => mult_143_n4199, B2 => B_SIG(10), C1 => 
                           mult_143_n4301, C2 => B_SIG(9), ZN => mult_143_n1815
                           );
   mult_143_U3846 : OAI21_X1 port map( B1 => mult_143_n6630, B2 => 
                           mult_143_n4467, A => mult_143_n1911, ZN => 
                           mult_143_n904);
   mult_143_U4163 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(3), B1 => 
                           mult_143_n4468, B2 => B_SIG(2), C1 => mult_143_n4468
                           , C2 => B_SIG(1), ZN => mult_143_n1911);
   mult_143_U3440 : AOI22_X1 port map( A1 => n3788, A2 => n3771, B1 => n3789, 
                           B2 => n3762, ZN => mult_143_n5852);
   mult_143_U3437 : AOI22_X1 port map( A1 => n3787, A2 => n3771, B1 => n3788, 
                           B2 => n3762, ZN => mult_143_n5849);
   mult_143_U2429 : XNOR2_X1 port map( A => mult_143_n4802, B => mult_143_n4803
                           , ZN => SIG_in(7));
   mult_143_U2434 : AOI21_X1 port map( B1 => n4724, B2 => n963, A => 
                           mult_143_n6501, ZN => mult_143_n4803);
   mult_143_U2435 : NOR2_X1 port map( A1 => n4709, A2 => n951, ZN => 
                           mult_143_n4802);
   mult_143_U2426 : XNOR2_X1 port map( A => mult_143_n4800, B => n2710, ZN => 
                           SIG_in(8));
   mult_143_U3428 : AOI22_X1 port map( A1 => n4695, A2 => n3821, B1 => n3784, 
                           B2 => n3771, ZN => mult_143_n5840);
   mult_143_U3434 : AOI22_X1 port map( A1 => n3787, A2 => n3821, B1 => n3786, 
                           B2 => n3771, ZN => mult_143_n5846);
   mult_143_U3708 : AOI22_X1 port map( A1 => n3787, A2 => n3540, B1 => n3810, 
                           B2 => n3789, ZN => mult_143_n6065);
   mult_143_U4541 : OAI21_X1 port map( B1 => mult_143_n2798, B2 => 
                           mult_143_n4467, A => mult_143_n1907, ZN => 
                           mult_143_n1536);
   mult_143_U4253 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(7), B1 => 
                           mult_143_n4468, B2 => B_SIG(6), C1 => mult_143_n4468
                           , C2 => B_SIG(5), ZN => mult_143_n1907);
   mult_143_U2999 : AOI22_X1 port map( A1 => n3792, A2 => n3791, B1 => n3769, 
                           B2 => n3768, ZN => mult_143_n2772);
   mult_143_U2424 : NOR2_X1 port map( A1 => n4860, A2 => mult_143_n2868, ZN => 
                           mult_143_n4799);
   mult_143_U2425 : OAI21_X1 port map( B1 => mult_143_n6517, B2 => 
                           mult_143_n4800, A => mult_143_n6516, ZN => 
                           mult_143_n4798);
   mult_143_U2427 : AOI21_X1 port map( B1 => n2603, B2 => n963, A => 
                           mult_143_n4801, ZN => mult_143_n4800);
   mult_143_U2428 : OAI21_X1 port map( B1 => mult_143_n412, B2 => n4709, A => 
                           mult_143_n4348, ZN => mult_143_n4801);
   mult_143_U3931 : AOI222_X1 port map( A1 => n1026, A2 => mult_143_n4468, B1 
                           => n1031, B2 => mult_143_n4468, C1 => mult_143_n3228
                           , C2 => B_SIG(23), ZN => mult_143_n2334);
   mult_143_U2734 : AOI222_X1 port map( A1 => n4634, A2 => n2780, B1 => n4634, 
                           B2 => mult_143_n1897, C1 => n2780, C2 => 
                           mult_143_n1897, ZN => mult_143_n650);
   mult_143_U3556 : AOI22_X1 port map( A1 => n4871, A2 => n3537, B1 => n3823, 
                           B2 => n4765, ZN => mult_143_n5958);
   mult_143_U2747 : AOI222_X1 port map( A1 => n3795, A2 => n2780, B1 => n3795, 
                           B2 => mult_143_n1892, C1 => n2780, C2 => 
                           mult_143_n1892, ZN => mult_143_n581);
   mult_143_U4591 : OAI21_X1 port map( B1 => mult_143_n2919, B2 => 
                           mult_143_n4467, A => mult_143_n1906, ZN => n993);
   mult_143_U3710 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(8), B1 => 
                           mult_143_n4468, B2 => B_SIG(7), C1 => mult_143_n4468
                           , C2 => B_SIG(6), ZN => mult_143_n1906);
   mult_143_U2701 : AOI22_X1 port map( A1 => n3793, A2 => mult_143_n1528, B1 =>
                           n667, B2 => n3803, ZN => mult_143_n5068);
   mult_143_U3497 : AOI22_X1 port map( A1 => B_SIG(19), A2 => n1026, B1 => 
                           B_SIG(17), B2 => mult_143_n3228, ZN => 
                           mult_143_n5901);
   mult_143_U3503 : AOI22_X1 port map( A1 => n3788, A2 => n3808, B1 => n3786, 
                           B2 => n3536, ZN => mult_143_n5907);
   mult_143_U2438 : XNOR2_X1 port map( A => mult_143_n4805, B => mult_143_n4806
                           , ZN => SIG_in(4));
   mult_143_U2439 : NAND2_X1 port map( A1 => mult_143_n4359, A2 => n4731, ZN =>
                           mult_143_n4806);
   mult_143_U2687 : AOI22_X1 port map( A1 => n3516, A2 => n1552, B1 => 
                           mult_143_n1900, B2 => n3824, ZN => mult_143_n5059);
   mult_143_U3553 : AOI22_X1 port map( A1 => B_SIG(20), A2 => mult_143_n36, B1 
                           => B_SIG(22), B2 => n755, ZN => mult_143_n5955);
   mult_143_U3684 : AOI21_X1 port map( B1 => n778, B2 => B_SIG(4), A => 
                           mult_143_n6049, ZN => mult_143_n6048);
   mult_143_U3685 : OAI21_X1 port map( B1 => mult_143_n4842, B2 => 
                           mult_143_n6629, A => mult_143_n6050, ZN => 
                           mult_143_n6049);
   mult_143_U3766 : AOI21_X1 port map( B1 => B_SIG(22), B2 => B_SIG(21), A => 
                           mult_143_n6104, ZN => mult_143_n6103);
   mult_143_U3506 : AOI22_X1 port map( A1 => n3787, A2 => n3536, B1 => n3789, 
                           B2 => n3808, ZN => mult_143_n5910);
   mult_143_U3509 : AOI22_X1 port map( A1 => n4871, A2 => n3536, B1 => n4765, 
                           B2 => n3808, ZN => mult_143_n5913);
   mult_143_U2732 : AOI22_X1 port map( A1 => n3810, A2 => n4765, B1 => n4871, 
                           B2 => n3540, ZN => mult_143_n5094);
   mult_143_U2436 : XNOR2_X1 port map( A => n2601, B => mult_143_n4804, ZN => 
                           SIG_in(5));
   mult_143_U2437 : AOI21_X1 port map( B1 => mult_143_n4359, B2 => 
                           mult_143_n4805, A => mult_143_n6510, ZN => 
                           mult_143_n4804);
   mult_143_U2440 : OAI21_X1 port map( B1 => mult_143_n6496, B2 => 
                           mult_143_n6491, A => mult_143_n6490, ZN => 
                           mult_143_n4805);
   mult_143_U2706 : AOI22_X1 port map( A1 => n3810, A2 => n3788, B1 => n3540, 
                           B2 => n3786, ZN => mult_143_n5071);
   mult_143_U2708 : AOI22_X1 port map( A1 => n1551, A2 => n3692, B1 => n4601, 
                           B2 => mult_143_n1898, ZN => mult_143_n671);
   mult_143_U2710 : AOI22_X1 port map( A1 => A_SIG(8), A2 => n1828, B1 => 
                           mult_143_n1818, B2 => n1782, ZN => mult_143_n5074);
   mult_143_U3623 : AOI222_X1 port map( A1 => mult_143_n4325, A2 => B_SIG(8), 
                           B1 => mult_143_n4206, B2 => B_SIG(7), C1 => 
                           mult_143_n4307, C2 => B_SIG(6), ZN => mult_143_n1818
                           );
   mult_143_U3542 : AOI222_X1 port map( A1 => mult_143_n4327, A2 => B_SIG(10), 
                           B1 => mult_143_n4208, B2 => B_SIG(9), C1 => 
                           mult_143_n4309, C2 => B_SIG(8), ZN => mult_143_n1816
                           );
   mult_143_U3777 : NOR2_X1 port map( A1 => B_SIG(21), A2 => B_SIG(22), ZN => 
                           mult_143_n6104);
   mult_143_U2745 : XNOR2_X1 port map( A => n3795, B => mult_143_n5111, ZN => 
                           n975);
   mult_143_U2746 : AOI22_X1 port map( A1 => mult_143_n1521, A2 => n4760, B1 =>
                           n2780, B2 => mult_143_n1892, ZN => mult_143_n5111);
   mult_143_U2655 : AOI22_X1 port map( A1 => n3791, A2 => n1550, B1 => 
                           mult_143_n1902, B2 => mult_143_n6367, ZN => 
                           mult_143_n744);
   mult_143_U2607 : AOI22_X1 port map( A1 => n3791, A2 => n3589, B1 => n4579, 
                           B2 => n4670, ZN => mult_143_n4985);
   mult_143_U4240 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => 
                           mult_143_n4467, A => mult_143_n1905, ZN => n1549);
   mult_143_U4124 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(9), B1 => 
                           mult_143_n4468, B2 => B_SIG(8), C1 => mult_143_n4468
                           , C2 => B_SIG(7), ZN => mult_143_n1905);
   mult_143_U3564 : OAI21_X1 port map( B1 => mult_143_n6627, B2 => 
                           mult_143_n4467, A => mult_143_n1904, ZN => n1548);
   mult_143_U4125 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(10), B1 => 
                           mult_143_n4468, B2 => B_SIG(9), C1 => mult_143_n4468
                           , C2 => B_SIG(8), ZN => mult_143_n1904);
   mult_143_U3547 : AOI22_X1 port map( A1 => n4688, A2 => n3823, B1 => n3784, 
                           B2 => n3537, ZN => mult_143_n5949);
   mult_143_U3500 : AOI22_X1 port map( A1 => n3787, A2 => n3808, B1 => n3536, 
                           B2 => n3785, ZN => mult_143_n5904);
   mult_143_U3605 : AOI22_X1 port map( A1 => n4871, A2 => n3805, B1 => n3786, 
                           B2 => n3539, ZN => n1498);
   mult_143_U2682 : AOI22_X1 port map( A1 => n3810, A2 => n4688, B1 => n3540, 
                           B2 => n3784, ZN => mult_143_n5054);
   mult_143_U3679 : AOI22_X1 port map( A1 => n4871, A2 => n3533, B1 => n3825, 
                           B2 => n4765, ZN => mult_143_n6045);
   mult_143_U3688 : AOI21_X1 port map( B1 => n1027, B2 => B_SIG(4), A => 
                           mult_143_n6052, ZN => mult_143_n6051);
   mult_143_U3689 : OAI21_X1 port map( B1 => n1068, B2 => mult_143_n4842, A => 
                           mult_143_n6053, ZN => mult_143_n6052);
   mult_143_U3385 : AOI21_X1 port map( B1 => B_SIG(6), B2 => mult_143_n2, A => 
                           mult_143_n5800, ZN => mult_143_n5799);
   mult_143_U3386 : OAI21_X1 port map( B1 => mult_143_n5124, B2 => 
                           mult_143_n2800, A => mult_143_n5801, ZN => 
                           mult_143_n5800);
   mult_143_U3387 : AOI22_X1 port map( A1 => B_SIG(5), A2 => mult_143_n3245, B1
                           => B_SIG(4), B2 => n1030, ZN => mult_143_n5801);
   mult_143_U3518 : AOI21_X1 port map( B1 => B_SIG(5), B2 => n1023, A => 
                           mult_143_n5921, ZN => mult_143_n5920);
   mult_143_U3519 : OAI21_X1 port map( B1 => mult_143_n4848, B2 => 
                           mult_143_n2800, A => mult_143_n5922, ZN => 
                           mult_143_n5921);
   mult_143_U3454 : AOI221_X1 port map( B1 => B_SIG(3), B2 => n1031, C1 => 
                           B_SIG(2), C2 => mult_143_n3228, A => mult_143_n5861,
                           ZN => mult_143_n5860);
   mult_143_U3455 : OAI22_X1 port map( A1 => n2977, A2 => n1053, B1 => 
                           mult_143_n5859, B2 => mult_143_n6629, ZN => 
                           mult_143_n5861);
   mult_143_U3513 : AOI221_X1 port map( B1 => n1023, B2 => B_SIG(3), C1 => 
                           B_SIG(2), C2 => mult_143_n36, A => mult_143_n5917, 
                           ZN => mult_143_n5916);
   mult_143_U3514 : OAI22_X1 port map( A1 => n2977, A2 => n976, B1 => 
                           mult_143_n4848, B2 => mult_143_n6629, ZN => 
                           mult_143_n5917);
   mult_143_U2822 : AOI22_X1 port map( A1 => n3789, A2 => n3798, B1 => n3807, 
                           B2 => n4765, ZN => mult_143_n5203);
   mult_143_U3758 : NAND2_X1 port map( A1 => B_SIG(19), A2 => n851, ZN => 
                           mult_143_n6096);
   mult_143_U3038 : XNOR2_X1 port map( A => mult_143_n5475, B => n2730, ZN => 
                           mult_143_n5375);
   mult_143_U3039 : XNOR2_X1 port map( A => n4935, B => n3090, ZN => 
                           mult_143_n5475);
   mult_143_U2815 : AOI22_X1 port map( A1 => n778, A2 => B_SIG(10), B1 => 
                           mult_143_n84, B2 => B_SIG(8), ZN => mult_143_n5197);
   mult_143_U3391 : AOI21_X1 port map( B1 => B_SIG(8), B2 => mult_143_n2, A => 
                           mult_143_n5806, ZN => mult_143_n5805);
   mult_143_U3392 : OAI21_X1 port map( B1 => mult_143_n2919, B2 => 
                           mult_143_n5124, A => mult_143_n5807, ZN => 
                           mult_143_n5806);
   mult_143_U3393 : AOI22_X1 port map( A1 => B_SIG(7), A2 => mult_143_n3245, B1
                           => B_SIG(6), B2 => n1030, ZN => mult_143_n5807);
   mult_143_U3599 : AOI22_X1 port map( A1 => n3786, A2 => n3805, B1 => n3767, 
                           B2 => n3785, ZN => mult_143_n5998);
   mult_143_U3521 : AOI21_X1 port map( B1 => B_SIG(7), B2 => n1023, A => 
                           mult_143_n5924, ZN => mult_143_n5923);
   mult_143_U3522 : OAI21_X1 port map( B1 => mult_143_n2919, B2 => 
                           mult_143_n4848, A => mult_143_n5925, ZN => 
                           mult_143_n5924);
   mult_143_U3523 : AOI22_X1 port map( A1 => B_SIG(6), A2 => mult_143_n36, B1 
                           => B_SIG(8), B2 => n755, ZN => mult_143_n5925);
   mult_143_U3465 : AOI21_X1 port map( B1 => B_SIG(7), B2 => n1031, A => 
                           mult_143_n5870, ZN => mult_143_n5869);
   mult_143_U3466 : OAI21_X1 port map( B1 => mult_143_n2919, B2 => 
                           mult_143_n5859, A => mult_143_n5871, ZN => 
                           mult_143_n5870);
   mult_143_U3467 : AOI22_X1 port map( A1 => B_SIG(6), A2 => mult_143_n3228, B1
                           => B_SIG(8), B2 => n1026, ZN => mult_143_n5871);
   mult_143_U3786 : OAI21_X1 port map( B1 => B_SIG(21), B2 => B_SIG(23), A => 
                           B_SIG(22), ZN => mult_143_n6123);
   mult_143_U2697 : AOI22_X1 port map( A1 => n3787, A2 => n3646, B1 => n3540, 
                           B2 => n3785, ZN => mult_143_n5065);
   mult_143_U3806 : AOI21_X1 port map( B1 => B_SIG(21), B2 => B_SIG(23), A => 
                           B_SIG(22), ZN => mult_143_n6122);
   mult_143_U2480 : AOI22_X1 port map( A1 => n4675, A2 => n3537, B1 => n4747, 
                           B2 => n3817, ZN => mult_143_n4858);
   mult_143_U3537 : NAND2_X1 port map( A1 => mult_143_n5940, A2 => n636, ZN => 
                           mult_143_n5938);
   mult_143_U2653 : AOI22_X1 port map( A1 => n778, A2 => B_SIG(17), B1 => 
                           mult_143_n84, B2 => B_SIG(15), ZN => mult_143_n5028)
                           ;
   mult_143_U3516 : AOI221_X1 port map( B1 => n755, B2 => B_SIG(5), C1 => 
                           B_SIG(3), C2 => mult_143_n36, A => mult_143_n5919, 
                           ZN => mult_143_n5918);
   mult_143_U3517 : OAI22_X1 port map( A1 => n1068, A2 => mult_143_n4848, B1 =>
                           n2977, B2 => n974, ZN => mult_143_n5919);
   mult_143_U3457 : AOI221_X1 port map( B1 => B_SIG(5), B2 => n1026, C1 => 
                           B_SIG(3), C2 => mult_143_n3228, A => mult_143_n5863,
                           ZN => mult_143_n5862);
   mult_143_U3458 : OAI22_X1 port map( A1 => n1068, A2 => mult_143_n5859, B1 =>
                           n2977, B2 => n980, ZN => mult_143_n5863);
   mult_143_U3560 : AOI221_X1 port map( B1 => B_SIG(5), B2 => n765, C1 => 
                           B_SIG(3), C2 => mult_143_n48, A => mult_143_n5962, 
                           ZN => mult_143_n5961);
   mult_143_U3561 : OAI22_X1 port map( A1 => n1068, A2 => mult_143_n4828, B1 =>
                           n2977, B2 => n1052, ZN => mult_143_n5962);
   mult_143_U3751 : AOI21_X1 port map( B1 => B_SIG(17), B2 => B_SIG(18), A => 
                           mult_143_n6003, ZN => mult_143_n6089);
   mult_143_U3696 : AOI21_X1 port map( B1 => n1027, B2 => B_SIG(7), A => 
                           mult_143_n6058, ZN => mult_143_n6057);
   mult_143_U3697 : OAI21_X1 port map( B1 => mult_143_n2919, B2 => 
                           mult_143_n4842, A => mult_143_n6059, ZN => 
                           mult_143_n6058);
   mult_143_U3698 : AOI22_X1 port map( A1 => n778, A2 => B_SIG(8), B1 => 
                           mult_143_n84, B2 => B_SIG(6), ZN => mult_143_n6059);
   mult_143_U3615 : AOI21_X1 port map( B1 => B_SIG(7), B2 => n774, A => 
                           mult_143_n6013, ZN => mult_143_n6012);
   mult_143_U3616 : OAI21_X1 port map( B1 => mult_143_n2919, B2 => 
                           mult_143_n4824, A => mult_143_n6014, ZN => 
                           mult_143_n6013);
   mult_143_U3617 : AOI22_X1 port map( A1 => B_SIG(6), A2 => mult_143_n72, B1 
                           => B_SIG(8), B2 => n772, ZN => mult_143_n6014);
   mult_143_U3756 : AOI22_X1 port map( A1 => n4714, A2 => n3772, B1 => n4688, 
                           B2 => n3531, ZN => mult_143_n6093);
   mult_143_U2519 : AOI22_X1 port map( A1 => n4871, A2 => n3823, B1 => n4688, 
                           B2 => n3799, ZN => mult_143_n4902);
   mult_143_U2545 : AOI22_X1 port map( A1 => n3810, A2 => n3827, B1 => n3540, 
                           B2 => n3777, ZN => mult_143_n4924);
   mult_143_U2769 : NAND2_X1 port map( A1 => mult_143_n5132, A2 => 
                           mult_143_n5133, ZN => n1715);
   mult_143_U2771 : AOI21_X1 port map( B1 => B_SIG(5), B2 => mult_143_n2, A => 
                           mult_143_n5135, ZN => mult_143_n5134);
   mult_143_U2772 : OAI21_X1 port map( B1 => n1068, B2 => mult_143_n5124, A => 
                           mult_143_n5136, ZN => mult_143_n5135);
   mult_143_U2773 : AOI22_X1 port map( A1 => B_SIG(3), A2 => n1030, B1 => 
                           B_SIG(4), B2 => mult_143_n3245, ZN => mult_143_n5136
                           );
   mult_143_U3816 : OAI22_X1 port map( A1 => n910, A2 => n1053, B1 => 
                           mult_143_n5859, B2 => mult_143_n3094, ZN => 
                           mult_143_n6134);
   mult_143_U3404 : AOI21_X1 port map( B1 => B_SIG(12), B2 => mult_143_n2, A =>
                           mult_143_n5818, ZN => mult_143_n5817);
   mult_143_U3405 : OAI21_X1 port map( B1 => mult_143_n6626, B2 => 
                           mult_143_n5124, A => mult_143_n5819, ZN => 
                           mult_143_n5818);
   mult_143_U3406 : AOI22_X1 port map( A1 => B_SIG(10), A2 => n1030, B1 => 
                           B_SIG(11), B2 => mult_143_n3245, ZN => 
                           mult_143_n5819);
   mult_143_U3462 : AOI21_X1 port map( B1 => B_SIG(6), B2 => n1031, A => 
                           mult_143_n5867, ZN => mult_143_n5866);
   mult_143_U3463 : OAI21_X1 port map( B1 => mult_143_n2798, B2 => 
                           mult_143_n5859, A => mult_143_n5868, ZN => 
                           mult_143_n5867);
   mult_143_U3464 : AOI22_X1 port map( A1 => B_SIG(5), A2 => mult_143_n3228, B1
                           => B_SIG(7), B2 => n1026, ZN => mult_143_n5868);
   mult_143_U3388 : AOI21_X1 port map( B1 => B_SIG(7), B2 => mult_143_n2, A => 
                           mult_143_n5803, ZN => mult_143_n5802);
   mult_143_U3389 : OAI21_X1 port map( B1 => mult_143_n2798, B2 => 
                           mult_143_n5124, A => mult_143_n5804, ZN => 
                           mult_143_n5803);
   mult_143_U3390 : AOI22_X1 port map( A1 => B_SIG(5), A2 => n1030, B1 => 
                           B_SIG(6), B2 => mult_143_n3245, ZN => mult_143_n5804
                           );
   mult_143_U3461 : OAI22_X1 port map( A1 => n895, A2 => n1053, B1 => 
                           mult_143_n5859, B2 => mult_143_n2800, ZN => 
                           mult_143_n5865);
   mult_143_U2508 : AOI22_X1 port map( A1 => mult_143_n74, A2 => B_SIG(9), B1 
                           => mult_143_n84, B2 => B_SIG(7), ZN => 
                           mult_143_n4888);
   mult_143_U3581 : AOI22_X1 port map( A1 => B_SIG(18), A2 => n787, B1 => 
                           B_SIG(17), B2 => mult_143_n48, ZN => mult_143_n5982)
                           ;
   mult_143_U3611 : AOI21_X1 port map( B1 => B_SIG(6), B2 => n774, A => 
                           mult_143_n6010, ZN => mult_143_n6009);
   mult_143_U3612 : OAI21_X1 port map( B1 => mult_143_n2798, B2 => 
                           mult_143_n4824, A => mult_143_n6011, ZN => 
                           mult_143_n6010);
   mult_143_U3613 : AOI22_X1 port map( A1 => B_SIG(5), A2 => mult_143_n72, B1 
                           => B_SIG(7), B2 => n772, ZN => mult_143_n6011);
   mult_143_U3692 : AOI21_X1 port map( B1 => n1027, B2 => B_SIG(6), A => 
                           mult_143_n6055, ZN => mult_143_n6054);
   mult_143_U3693 : OAI21_X1 port map( B1 => mult_143_n2798, B2 => 
                           mult_143_n4842, A => mult_143_n6056, ZN => 
                           mult_143_n6055);
   mult_143_U3694 : AOI22_X1 port map( A1 => n778, A2 => B_SIG(7), B1 => 
                           mult_143_n84, B2 => B_SIG(5), ZN => mult_143_n6056);
   mult_143_U3674 : AOI21_X1 port map( B1 => B_SIG(20), B2 => B_SIG(19), A => 
                           mult_143_n6042, ZN => mult_143_n6041);
   mult_143_U3675 : NOR2_X1 port map( A1 => B_SIG(20), A2 => B_SIG(19), ZN => 
                           mult_143_n6042);
   mult_143_U3725 : OAI21_X1 port map( B1 => n1068, B2 => mult_143_n4891, A => 
                           mult_143_n6073, ZN => mult_143_n6072);
   mult_143_U3726 : AOI22_X1 port map( A1 => B_SIG(5), A2 => n2598, B1 => 
                           B_SIG(3), B2 => mult_143_n96, ZN => mult_143_n6073);
   mult_143_U3721 : OAI21_X1 port map( B1 => mult_143_n4891, B2 => 
                           mult_143_n6629, A => mult_143_n6070, ZN => 
                           mult_143_n6069);
   mult_143_U3722 : AOI22_X1 port map( A1 => B_SIG(3), A2 => n799, B1 => 
                           B_SIG(2), B2 => mult_143_n96, ZN => mult_143_n6070);
   mult_143_U3042 : NAND2_X1 port map( A1 => mult_143_n5484, A2 => 
                           mult_143_n5485, ZN => n954);
   mult_143_U3055 : XNOR2_X1 port map( A => n3498, B => n3750, ZN => 
                           mult_143_n5495);
   mult_143_U3056 : AOI222_X1 port map( A1 => n3493, A2 => n1575, B1 => n3493, 
                           B2 => n3709, C1 => n1575, C2 => n3709, ZN => 
                           mult_143_n5484);
   mult_143_U3742 : NOR2_X1 port map( A1 => B_SIG(15), A2 => B_SIG(16), ZN => 
                           mult_143_n6085);
   mult_143_U2941 : AOI222_X1 port map( A1 => n2723, A2 => mult_143_n5274, B1 
                           => n2723, B2 => mult_143_n5273, C1 => mult_143_n5274
                           , C2 => mult_143_n5273, ZN => mult_143_n5265);
   mult_143_U3585 : AOI22_X1 port map( A1 => n3787, A2 => n3538, B1 => n3788, 
                           B2 => n3807, ZN => mult_143_n5985);
   mult_143_U2819 : AOI22_X1 port map( A1 => n3788, A2 => n3767, B1 => n3789, 
                           B2 => n3805, ZN => mult_143_n5200);
   mult_143_U2470 : AOI22_X1 port map( A1 => n1027, A2 => B_SIG(2), B1 => 
                           mult_143_n84, B2 => B_SIG(1), ZN => mult_143_n4843);
   mult_143_U3822 : NAND2_X1 port map( A1 => mult_143_n6135, A2 => 
                           mult_143_n6136, ZN => mult_143_n6138);
   mult_143_U3480 : AOI21_X1 port map( B1 => B_SIG(13), B2 => n1031, A => 
                           mult_143_n5885, ZN => mult_143_n5884);
   mult_143_U3481 : OAI21_X1 port map( B1 => mult_143_n3443, B2 => 
                           mult_143_n5859, A => mult_143_n5886, ZN => 
                           mult_143_n5885);
   mult_143_U3482 : AOI22_X1 port map( A1 => B_SIG(12), A2 => mult_143_n3228, 
                           B1 => B_SIG(14), B2 => n1026, ZN => mult_143_n5886);
   mult_143_U3411 : AOI21_X1 port map( B1 => B_SIG(14), B2 => mult_143_n2, A =>
                           mult_143_n5824, ZN => mult_143_n5823);
   mult_143_U3412 : OAI21_X1 port map( B1 => mult_143_n3443, B2 => 
                           mult_143_n5124, A => mult_143_n5825, ZN => 
                           mult_143_n5824);
   mult_143_U3413 : AOI22_X1 port map( A1 => B_SIG(13), A2 => mult_143_n3245, 
                           B1 => B_SIG(12), B2 => n1030, ZN => mult_143_n5825);
   mult_143_U3150 : XNOR2_X1 port map( A => mult_143_n5605, B => n3057, ZN => 
                           mult_143_n5587);
   mult_143_U3151 : XNOR2_X1 port map( A => n2874, B => n2829, ZN => 
                           mult_143_n5605);
   mult_143_U3877 : AOI22_X1 port map( A1 => B_SIG(9), A2 => n755, B1 => 
                           B_SIG(8), B2 => n1023, ZN => mult_143_n6194);
   mult_143_U2475 : AOI22_X1 port map( A1 => B_SIG(15), A2 => n1023, B1 => 
                           B_SIG(16), B2 => n755, ZN => mult_143_n4849);
   mult_143_U3078 : NAND2_X1 port map( A1 => mult_143_n5532, A2 => 
                           mult_143_n5533, ZN => n945);
   mult_143_U3353 : OAI21_X1 port map( B1 => n712, B2 => n3760, A => 
                           mult_143_n5775, ZN => mult_143_n218);
   mult_143_U3354 : OAI21_X1 port map( B1 => n1711, B2 => n712, A => n3760, ZN 
                           => mult_143_n5775);
   mult_143_U3355 : XNOR2_X1 port map( A => mult_143_n5776, B => mult_143_n5777
                           , ZN => n1714);
   mult_143_U3356 : XNOR2_X1 port map( A => mult_143_n5778, B => mult_143_n5779
                           , ZN => mult_143_n5777);
   mult_143_U3357 : AOI222_X1 port map( A1 => mult_143_n5782, A2 => n4634, B1 
                           => mult_143_n5782, B2 => n2617, C1 => n4634, C2 => 
                           n2617, ZN => mult_143_n5781);
   mult_143_U3358 : XNOR2_X1 port map( A => mult_143_n5783, B => mult_143_n5784
                           , ZN => mult_143_n5780);
   mult_143_U3359 : XNOR2_X1 port map( A => mult_143_n6309, B => n4752, ZN => 
                           mult_143_n5784);
   mult_143_U3362 : OAI21_X1 port map( B1 => n1711, B2 => n3515, A => n1712, ZN
                           => mult_143_n5787);
   mult_143_U3450 : XNOR2_X1 port map( A => A_SIG(5), B => mult_143_n5857, ZN 
                           => n1713);
   mult_143_U3451 : AOI221_X1 port map( B1 => B_SIG(3), B2 => n1026, C1 => 
                           B_SIG(1), C2 => mult_143_n3228, A => mult_143_n5858,
                           ZN => mult_143_n5857);
   mult_143_U3452 : OAI22_X1 port map( A1 => mult_143_n6630, A2 => 
                           mult_143_n5859, B1 => n910, B2 => n980, ZN => 
                           mult_143_n5858);
   mult_143_U3080 : XNOR2_X1 port map( A => mult_143_n5534, B => n3515, ZN => 
                           mult_143_n5533);
   mult_143_U3364 : AOI222_X1 port map( A1 => mult_143_n5542, A2 => 
                           mult_143_n5543, B1 => mult_143_n5542, B2 => 
                           mult_143_n5540, C1 => mult_143_n5543, C2 => 
                           mult_143_n5540, ZN => n1494);
   mult_143_U3081 : NOR2_X1 port map( A1 => n1711, A2 => n2762, ZN => 
                           mult_143_n5534);
   mult_143_U3363 : NAND2_X1 port map( A1 => n3757, A2 => n3758, ZN => n1712);
   mult_143_U3374 : NOR2_X1 port map( A1 => n3758, A2 => n3757, ZN => n1711);
   mult_143_U3375 : XNOR2_X1 port map( A => mult_143_n5782, B => mult_143_n5794
                           , ZN => mult_143_n5789);
   mult_143_U3377 : XNOR2_X1 port map( A => n2633, B => n2751, ZN => 
                           mult_143_n5782);
   mult_143_U3378 : XNOR2_X1 port map( A => mult_143_n5786, B => mult_143_n5796
                           , ZN => mult_143_n5788);
   mult_143_U3384 : AOI222_X1 port map( A1 => mult_143_n1893, A2 => n2630, B1 
                           => mult_143_n1893, B2 => n2733, C1 => n2630, C2 => 
                           n2733, ZN => mult_143_n5786);
   mult_143_U3082 : AOI222_X1 port map( A1 => n3512, A2 => n3747, B1 => n3512, 
                           B2 => n3700, C1 => n3747, C2 => n3700, ZN => 
                           mult_143_n5532);
   mult_143_U2650 : AOI22_X1 port map( A1 => n3789, A2 => n3767, B1 => n4765, 
                           B2 => n3805, ZN => mult_143_n5025);
   mult_143_U3534 : OAI21_X1 port map( B1 => n3673, B2 => n3667, A => 
                           mult_143_n5937, ZN => mult_143_n5936);
   mult_143_U3535 : AOI22_X1 port map( A1 => n3537, A2 => n3779, B1 => n3781, 
                           B2 => n3823, ZN => mult_143_n5937);
   mult_143_U3342 : XNOR2_X1 port map( A => n4652, B => n2664, ZN => 
                           mult_143_n5768);
   mult_143_U2685 : AOI22_X1 port map( A1 => B_SIG(21), A2 => n774, B1 => n772,
                           B2 => B_SIG(22), ZN => mult_143_n5057);
   mult_143_U3468 : AOI21_X1 port map( B1 => B_SIG(8), B2 => n1031, A => 
                           mult_143_n5873, ZN => mult_143_n5872);
   mult_143_U3469 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => 
                           mult_143_n5859, A => mult_143_n5874, ZN => 
                           mult_143_n5873);
   mult_143_U3470 : AOI22_X1 port map( A1 => B_SIG(7), A2 => mult_143_n3228, B1
                           => B_SIG(9), B2 => n1026, ZN => mult_143_n5874);
   mult_143_U2668 : AOI22_X1 port map( A1 => n3788, A2 => n3825, B1 => n4688, 
                           B2 => n3533, ZN => mult_143_n5041);
   mult_143_U3395 : AOI21_X1 port map( B1 => B_SIG(9), B2 => mult_143_n2, A => 
                           mult_143_n5809, ZN => mult_143_n5808);
   mult_143_U3396 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => 
                           mult_143_n5124, A => mult_143_n5810, ZN => 
                           mult_143_n5809);
   mult_143_U3397 : AOI22_X1 port map( A1 => B_SIG(7), A2 => n1030, B1 => 
                           B_SIG(8), B2 => mult_143_n3245, ZN => mult_143_n5810
                           );
   mult_143_U2636 : AOI22_X1 port map( A1 => B_SIG(18), A2 => n774, B1 => 
                           B_SIG(17), B2 => mult_143_n72, ZN => mult_143_n5012)
                           ;
   mult_143_U2631 : AOI21_X1 port map( B1 => n3778, B2 => n3531, A => 
                           mult_143_n5008, ZN => mult_143_n5007);
   mult_143_U2594 : AOI22_X1 port map( A1 => B_SIG(15), A2 => mult_143_n72, B1 
                           => B_SIG(16), B2 => n774, ZN => mult_143_n4971);
   mult_143_U3818 : AOI21_X1 port map( B1 => B_SIG(3), B2 => n755, A => 
                           mult_143_n6140, ZN => mult_143_n6139);
   mult_143_U3819 : OAI21_X1 port map( B1 => mult_143_n6630, B2 => 
                           mult_143_n4848, A => mult_143_n6141, ZN => 
                           mult_143_n6140);
   mult_143_U3035 : AOI222_X1 port map( A1 => n966, A2 => n2888, B1 => n966, B2
                           => n4685, C1 => n2888, C2 => n4685, ZN => 
                           mult_143_n5372);
   mult_143_U3069 : AND2_X1 port map( A1 => n3511, A2 => n4637, ZN => 
                           mult_143_n5516);
   mult_143_U3303 : XNOR2_X1 port map( A => mult_143_n5738, B => n2666, ZN => 
                           mult_143_n5723);
   mult_143_U3304 : XNOR2_X1 port map( A => n2624, B => n4754, ZN => 
                           mult_143_n5738);
   mult_143_U3173 : XNOR2_X1 port map( A => mult_143_n5624, B => mult_143_n5617
                           , ZN => n1710);
   mult_143_U3175 : XNOR2_X1 port map( A => n4874, B => mult_143_n5616, ZN => 
                           mult_143_n5624);
   mult_143_U3011 : AOI22_X1 port map( A1 => n4695, A2 => n3825, B1 => n3783, 
                           B2 => n3533, ZN => mult_143_n5444);
   mult_143_U2444 : XNOR2_X1 port map( A => mult_143_n4810, B => mult_143_n4811
                           , ZN => mult_143_n994);
   mult_143_U2781 : XNOR2_X1 port map( A => n3513, B => n3752, ZN => 
                           mult_143_n5145);
   mult_143_U2782 : AOI222_X1 port map( A1 => n3738, A2 => n3500, B1 => n3738, 
                           B2 => n3754, C1 => n3500, C2 => n3754, ZN => 
                           mult_143_n5143);
   mult_143_U2988 : XNOR2_X1 port map( A => mult_143_n5415, B => mult_143_n5178
                           , ZN => n1708);
   mult_143_U2990 : XNOR2_X1 port map( A => n4671, B => n2610, ZN => 
                           mult_143_n5415);
   mult_143_U2859 : XNOR2_X1 port map( A => mult_143_n5273, B => mult_143_n5274
                           , ZN => mult_143_n5272);
   mult_143_U2945 : NOR2_X1 port map( A1 => mult_143_n5367, A2 => 
                           mult_143_n5368, ZN => mult_143_n5274);
   mult_143_U2946 : NOR2_X1 port map( A1 => n1757, A2 => n2938, ZN => 
                           mult_143_n5368);
   mult_143_U2947 : AOI21_X1 port map( B1 => n2938, B2 => n1757, A => n3636, ZN
                           => mult_143_n5367);
   mult_143_U2604 : AOI22_X1 port map( A1 => n3786, A2 => n3767, B1 => n3785, 
                           B2 => n4664, ZN => mult_143_n4981);
   mult_143_U2566 : AOI22_X1 port map( A1 => n3788, A2 => n3802, B1 => n3786, 
                           B2 => n3798, ZN => mult_143_n4946);
   mult_143_U3240 : XNOR2_X1 port map( A => mult_143_n6592, B => mult_143_n5673
                           , ZN => mult_143_n5648);
   mult_143_U2465 : AOI22_X1 port map( A1 => B_SIG(9), A2 => n804, B1 => 
                           B_SIG(8), B2 => mult_143_n6621, ZN => mult_143_n4839
                           );
   mult_143_U3400 : AOI22_X1 port map( A1 => B_SIG(9), A2 => mult_143_n3245, B1
                           => B_SIG(8), B2 => n1030, ZN => mult_143_n5813);
   mult_143_U3471 : AOI21_X1 port map( B1 => B_SIG(9), B2 => n1031, A => 
                           mult_143_n5876, ZN => mult_143_n5875);
   mult_143_U3472 : OAI21_X1 port map( B1 => mult_143_n6627, B2 => 
                           mult_143_n5859, A => mult_143_n5877, ZN => 
                           mult_143_n5876);
   mult_143_U3473 : AOI22_X1 port map( A1 => B_SIG(10), A2 => n1026, B1 => 
                           B_SIG(8), B2 => mult_143_n3228, ZN => mult_143_n5877
                           );
   mult_143_U3524 : AOI21_X1 port map( B1 => B_SIG(9), B2 => n1023, A => 
                           mult_143_n5927, ZN => mult_143_n5926);
   mult_143_U3525 : OAI21_X1 port map( B1 => mult_143_n6627, B2 => 
                           mult_143_n4848, A => mult_143_n5928, ZN => 
                           mult_143_n5927);
   mult_143_U3526 : AOI22_X1 port map( A1 => B_SIG(10), A2 => n755, B1 => 
                           B_SIG(8), B2 => mult_143_n36, ZN => mult_143_n5928);
   mult_143_U3562 : AOI21_X1 port map( B1 => B_SIG(10), B2 => n765, A => 
                           mult_143_n5964, ZN => mult_143_n5963);
   mult_143_U3563 : OAI21_X1 port map( B1 => mult_143_n6627, B2 => 
                           mult_143_n4828, A => mult_143_n5965, ZN => 
                           mult_143_n5964);
   mult_143_U3566 : AOI22_X1 port map( A1 => B_SIG(9), A2 => n787, B1 => 
                           B_SIG(8), B2 => mult_143_n48, ZN => mult_143_n5965);
   mult_143_U2933 : AOI222_X1 port map( A1 => mult_143_n5355, A2 => 
                           mult_143_n5354, B1 => mult_143_n5354, B2 => 
                           mult_143_n5356, C1 => mult_143_n5355, C2 => 
                           mult_143_n5356, ZN => mult_143_n5264);
   mult_143_U2938 : XNOR2_X1 port map( A => n4843, B => mult_143_n5361, ZN => 
                           mult_143_n5356);
   mult_143_U2939 : XNOR2_X1 port map( A => n4583, B => mult_143_n5362, ZN => 
                           mult_143_n5355);
   mult_143_U2940 : AOI222_X1 port map( A1 => n2728, A2 => n2621, B1 => n2728, 
                           B2 => mult_143_n5363, C1 => n2621, C2 => 
                           mult_143_n5363, ZN => mult_143_n5354);
   mult_143_U2942 : NOR2_X1 port map( A1 => mult_143_n5365, A2 => 
                           mult_143_n5366, ZN => mult_143_n5363);
   mult_143_U2943 : NOR2_X1 port map( A1 => n4615, A2 => n3634, ZN => 
                           mult_143_n5366);
   mult_143_U2944 : AOI21_X1 port map( B1 => n3634, B2 => n4615, A => n3621, ZN
                           => mult_143_n5365);
   mult_143_U2484 : AOI22_X1 port map( A1 => n3827, A2 => n3805, B1 => n3777, 
                           B2 => n4664, ZN => mult_143_n4861);
   mult_143_U3044 : AOI21_X1 port map( B1 => B_SIG(5), B2 => n1027, A => 
                           mult_143_n5487, ZN => mult_143_n5486);
   mult_143_U3045 : OAI21_X1 port map( B1 => mult_143_n4842, B2 => 
                           mult_143_n2800, A => mult_143_n5488, ZN => 
                           mult_143_n5487);
   mult_143_U3046 : AOI22_X1 port map( A1 => n778, A2 => B_SIG(6), B1 => 
                           mult_143_n84, B2 => B_SIG(4), ZN => mult_143_n5488);
   mult_143_U2787 : XNOR2_X1 port map( A => n4662, B => mult_143_n5161, ZN => 
                           mult_143_n5158);
   mult_143_U2788 : XNOR2_X1 port map( A => mult_143_n5163, B => mult_143_n5162
                           , ZN => n1707);
   mult_143_U2789 : XNOR2_X1 port map( A => n3106, B => mult_143_n5164, ZN => 
                           mult_143_n5162);
   mult_143_U2790 : AOI222_X1 port map( A1 => mult_143_n5165, A2 => n4888, B1 
                           => mult_143_n5165, B2 => n2796, C1 => n4888, C2 => 
                           n2796, ZN => n1493);
   mult_143_U3289 : XNOR2_X1 port map( A => mult_143_n5718, B => mult_143_n5717
                           , ZN => n1706);
   mult_143_U3290 : XNOR2_X1 port map( A => mult_143_n5719, B => mult_143_n5720
                           , ZN => mult_143_n5717);
   mult_143_U3227 : XNOR2_X1 port map( A => mult_143_n5666, B => mult_143_n6379
                           , ZN => mult_143_n5164);
   mult_143_U3417 : AOI21_X1 port map( B1 => n4747, B2 => n3801, A => 
                           mult_143_n5830, ZN => n1547);
   mult_143_U3418 : OAI21_X1 port map( B1 => n3655, B2 => n3659, A => n3530, ZN
                           => mult_143_n5830);
   mult_143_U3419 : AOI22_X1 port map( A1 => B_SIG(14), A2 => n1030, B1 => 
                           B_SIG(15), B2 => mult_143_n3245, ZN => 
                           mult_143_n5831);
   mult_143_U3488 : AOI22_X1 port map( A1 => n3781, A2 => n3536, B1 => n3783, 
                           B2 => n3808, ZN => mult_143_n5892);
   mult_143_U3576 : AOI21_X1 port map( B1 => n3783, B2 => n3802, A => 
                           mult_143_n5978, ZN => n1545);
   mult_143_U3577 : OAI21_X1 port map( B1 => n3655, B2 => n4734, A => n3529, ZN
                           => mult_143_n5978);
   mult_143_U3578 : AOI22_X1 port map( A1 => B_SIG(14), A2 => mult_143_n48, B1 
                           => B_SIG(15), B2 => n787, ZN => mult_143_n5979);
   mult_143_U2812 : AOI22_X1 port map( A1 => B_SIG(15), A2 => n804, B1 => 
                           B_SIG(16), B2 => n2599, ZN => mult_143_n5194);
   mult_143_U3057 : NAND2_X1 port map( A1 => mult_143_n5502, A2 => 
                           mult_143_n5503, ZN => n946);
   mult_143_U3059 : XNOR2_X1 port map( A => n3511, B => mult_143_n5504, ZN => 
                           mult_143_n5503);
   mult_143_U3060 : AOI22_X1 port map( A1 => n3746, A2 => n4637, B1 => n3699, 
                           B2 => n4639, ZN => mult_143_n5504);
   mult_143_U3061 : AOI222_X1 port map( A1 => n3498, A2 => n3750, B1 => n3498, 
                           B2 => n3591, C1 => n3750, C2 => n3591, ZN => 
                           mult_143_n5502);
   mult_143_U3063 : XNOR2_X1 port map( A => mult_143_n5509, B => mult_143_n5510
                           , ZN => n1705);
   mult_143_U3064 : XNOR2_X1 port map( A => mult_143_n5511, B => mult_143_n5512
                           , ZN => mult_143_n5509);
   mult_143_U3327 : AOI222_X1 port map( A1 => mult_143_n6346, A2 => n2627, B1 
                           => mult_143_n6346, B2 => n2667, C1 => n2627, C2 => 
                           n2667, ZN => mult_143_n5514);
   mult_143_U3728 : AOI21_X1 port map( B1 => B_SIG(9), B2 => n799, A => 
                           mult_143_n6075, ZN => mult_143_n6074);
   mult_143_U3729 : OAI21_X1 port map( B1 => mult_143_n6627, B2 => 
                           mult_143_n4891, A => mult_143_n6076, ZN => 
                           mult_143_n6075);
   mult_143_U3730 : AOI22_X1 port map( A1 => B_SIG(10), A2 => n2598, B1 => 
                           B_SIG(8), B2 => mult_143_n96, ZN => mult_143_n6076);
   mult_143_U3474 : AOI21_X1 port map( B1 => B_SIG(10), B2 => n1031, A => 
                           mult_143_n5879, ZN => mult_143_n5878);
   mult_143_U3476 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n1026, B1 => 
                           B_SIG(9), B2 => mult_143_n3228, ZN => mult_143_n5880
                           );
   mult_143_U3403 : AOI22_X1 port map( A1 => n3778, A2 => n3821, B1 => n3777, 
                           B2 => n4694, ZN => mult_143_n5816);
   mult_143_U2760 : OAI221_X1 port map( B1 => mult_143_n5118, B2 => 
                           mult_143_n5117, C1 => mult_143_n5122, C2 => A_SIG(2)
                           , A => mult_143_n5123, ZN => mult_143_n5121);
   mult_143_U2761 : NAND2_X1 port map( A1 => mult_143_n5122, A2 => A_SIG(2), ZN
                           => mult_143_n5123);
   mult_143_U2762 : OAI211_X1 port map( C1 => mult_143_n6630, C2 => 
                           mult_143_n5124, A => mult_143_n5125, B => 
                           mult_143_n5126, ZN => mult_143_n5122);
   mult_143_U2763 : NAND2_X1 port map( A1 => B_SIG(3), A2 => mult_143_n2, ZN =>
                           mult_143_n5126);
   mult_143_U2764 : AOI22_X1 port map( A1 => B_SIG(1), A2 => n1030, B1 => 
                           B_SIG(2), B2 => mult_143_n3245, ZN => mult_143_n5125
                           );
   mult_143_U2766 : AOI21_X1 port map( B1 => B_SIG(4), B2 => mult_143_n2, A => 
                           mult_143_n5130, ZN => mult_143_n5129);
   mult_143_U2767 : OAI21_X1 port map( B1 => mult_143_n5124, B2 => 
                           mult_143_n6629, A => mult_143_n5131, ZN => 
                           mult_143_n5130);
   mult_143_U2562 : AOI22_X1 port map( A1 => B_SIG(17), A2 => n804, B1 => 
                           B_SIG(16), B2 => mult_143_n6621, ZN => 
                           mult_143_n4943);
   mult_143_U3145 : XNOR2_X1 port map( A => mult_143_n5595, B => n2846, ZN => 
                           mult_143_n5576);
   mult_143_U3186 : XNOR2_X1 port map( A => n2668, B => n2767, ZN => 
                           mult_143_n5632);
   mult_143_U3420 : AOI21_X1 port map( B1 => B_SIG(17), B2 => mult_143_n2, A =>
                           mult_143_n5833, ZN => n1544);
   mult_143_U3422 : AOI22_X1 port map( A1 => B_SIG(15), A2 => n1030, B1 => 
                           B_SIG(16), B2 => mult_143_n3245, ZN => 
                           mult_143_n5834);
   mult_143_U3489 : AOI21_X1 port map( B1 => n4747, B2 => n3809, A => 
                           mult_143_n5894, ZN => mult_143_n5893);
   mult_143_U3491 : AOI22_X1 port map( A1 => n3784, A2 => n3808, B1 => n4675, 
                           B2 => n3536, ZN => mult_143_n5895);
   mult_143_U3963 : AOI222_X1 port map( A1 => n3722, A2 => n3725, B1 => n3722, 
                           B2 => n3520, C1 => n3725, C2 => n3520, ZN => 
                           mult_143_n1017);
   mult_143_U3527 : AOI21_X1 port map( B1 => B_SIG(10), B2 => n1023, A => 
                           mult_143_n5930, ZN => mult_143_n5929);
   mult_143_U3529 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n755, B1 => 
                           B_SIG(9), B2 => mult_143_n36, ZN => mult_143_n5931);
   mult_143_U3567 : AOI21_X1 port map( B1 => n3827, B2 => n3802, A => 
                           mult_143_n5967, ZN => mult_143_n5966);
   mult_143_U3860 : XNOR2_X1 port map( A => n649, B => mult_143_n6179, ZN => 
                           n1703);
   mult_143_U3861 : AOI221_X1 port map( B1 => n2599, B2 => B_SIG(3), C1 => 
                           B_SIG(1), C2 => mult_143_n6621, A => mult_143_n6180,
                           ZN => mult_143_n6179);
   mult_143_U3862 : OAI22_X1 port map( A1 => mult_143_n6630, A2 => 
                           mult_143_n4820, B1 => n910, B2 => n979, ZN => 
                           mult_143_n6180);
   mult_143_U3868 : OAI22_X1 port map( A1 => n910, A2 => n996, B1 => 
                           mult_143_n4820, B2 => n2817, ZN => mult_143_n6183);
   mult_143_U3594 : AOI21_X1 port map( B1 => n4747, B2 => n4665, A => 
                           mult_143_n5994, ZN => n1543);
   mult_143_U3596 : AOI22_X1 port map( A1 => n3784, A2 => n3805, B1 => n4675, 
                           B2 => n3539, ZN => mult_143_n5995);
   mult_143_U2830 : OAI21_X1 port map( B1 => n3746, B2 => n3699, A => 
                           mult_143_n5219, ZN => mult_143_n3073);
   mult_143_U2831 : AOI221_X1 port map( B1 => n4637, B2 => n3511, C1 => n4639, 
                           C2 => n3511, A => mult_143_n5221, ZN => 
                           mult_143_n5219);
   mult_143_U3068 : XNOR2_X1 port map( A => n3512, B => n3747, ZN => 
                           mult_143_n5517);
   mult_143_U3083 : XNOR2_X1 port map( A => mult_143_n5540, B => mult_143_n5541
                           , ZN => n1702);
   mult_143_U3373 : XNOR2_X1 port map( A => n2733, B => mult_143_n5793, ZN => 
                           mult_143_n5542);
   mult_143_U3365 : AOI222_X1 port map( A1 => mult_143_n6322, A2 => 
                           mult_143_n5527, B1 => mult_143_n6322, B2 => 
                           mult_143_n5525, C1 => mult_143_n5527, C2 => 
                           mult_143_n5525, ZN => mult_143_n5540);
   mult_143_U3084 : AOI222_X1 port map( A1 => mult_143_n5521, A2 => 
                           mult_143_n5523, B1 => mult_143_n5521, B2 => n2861, 
                           C1 => mult_143_n5523, C2 => n2861, ZN => n1491);
   mult_143_U3072 : NOR2_X1 port map( A1 => mult_143_n5528, A2 => 
                           mult_143_n5529, ZN => mult_143_n5505);
   mult_143_U3073 : NOR2_X1 port map( A1 => mult_143_n6582, A2 => 
                           mult_143_n6581, ZN => mult_143_n5529);
   mult_143_U3075 : XNOR2_X1 port map( A => mult_143_n5530, B => n3794, ZN => 
                           mult_143_n5508);
   mult_143_U3076 : XNOR2_X1 port map( A => n2631, B => n3625, ZN => 
                           mult_143_n5530);
   mult_143_U3077 : OAI222_X1 port map( A1 => n2692, A2 => n2714, B1 => 
                           mult_143_n5531, B2 => n2692, C1 => mult_143_n5531, 
                           C2 => n2714, ZN => mult_143_n5507);
   mult_143_U3368 : AOI21_X1 port map( B1 => n4760, B2 => n4632, A => 
                           mult_143_n5791, ZN => mult_143_n5527);
   mult_143_U3369 : AOI21_X1 port map( B1 => n2749, B2 => mult_143_n4490, A => 
                           n3056, ZN => mult_143_n5791);
   mult_143_U3366 : XNOR2_X1 port map( A => n3051, B => n2751, ZN => 
                           mult_143_n5525);
   mult_143_U3070 : XNOR2_X1 port map( A => mult_143_n5522, B => mult_143_n5521
                           , ZN => n1701);
   mult_143_U3086 : NOR2_X1 port map( A1 => mult_143_n5544, A2 => 
                           mult_143_n5545, ZN => mult_143_n5510);
   mult_143_U3087 : NOR2_X1 port map( A1 => n3054, A2 => n2732, ZN => 
                           mult_143_n5545);
   mult_143_U3088 : AOI21_X1 port map( B1 => n2732, B2 => n3054, A => 
                           mult_143_n1896, ZN => mult_143_n5544);
   mult_143_U3089 : XNOR2_X1 port map( A => n2731, B => mult_143_n1895, ZN => 
                           mult_143_n5512);
   mult_143_U3091 : XNOR2_X1 port map( A => n3056, B => mult_143_n5547, ZN => 
                           mult_143_n5511);
   mult_143_U3092 : AOI22_X1 port map( A1 => n2749, A2 => n4632, B1 => 
                           mult_143_n4490, B2 => n4760, ZN => mult_143_n5547);
   mult_143_U3093 : XNOR2_X1 port map( A => n2620, B => mult_143_n1523, ZN => 
                           mult_143_n5523);
   mult_143_U3100 : AOI222_X1 port map( A1 => n2631, A2 => n3625, B1 => n2631, 
                           B2 => n3794, C1 => n3625, C2 => n3794, ZN => 
                           mult_143_n5521);
   mult_143_U2503 : AOI22_X1 port map( A1 => n3779, A2 => n3539, B1 => n4736, 
                           B2 => n3805, ZN => mult_143_n4881);
   mult_143_U3660 : AOI21_X1 port map( B1 => n4675, B2 => n3819, A => 
                           mult_143_n6033, ZN => n1542);
   mult_143_U3661 : OAI21_X1 port map( B1 => n3655, B2 => n3596, A => n3528, ZN
                           => mult_143_n6033);
   mult_143_U3662 : AOI22_X1 port map( A1 => B_SIG(14), A2 => mult_143_n72, B1 
                           => B_SIG(16), B2 => n772, ZN => mult_143_n6034);
   mult_143_U3264 : AOI222_X1 port map( A1 => n3735, A2 => n4568, B1 => n3735, 
                           B2 => n1687, C1 => n4568, C2 => n1687, ZN => 
                           mult_143_n5697);
   mult_143_U2499 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n772, B1 => 
                           B_SIG(9), B2 => mult_143_n72, ZN => mult_143_n4878);
   mult_143_U3206 : XNOR2_X1 port map( A => mult_143_n5649, B => mult_143_n5650
                           , ZN => n1700);
   mult_143_U3207 : XNOR2_X1 port map( A => mult_143_n5651, B => mult_143_n5652
                           , ZN => mult_143_n5649);
   mult_143_U2931 : XNOR2_X1 port map( A => mult_143_n5353, B => mult_143_n6434
                           , ZN => mult_143_n5253);
   mult_143_U2932 : XNOR2_X1 port map( A => mult_143_n6432, B => n2803, ZN => 
                           mult_143_n5353);
   mult_143_U2366 : NAND2_X1 port map( A1 => n2764, A2 => n945, ZN => 
                           mult_143_n4756);
   mult_143_U2386 : OAI21_X1 port map( B1 => n726, B2 => mult_143_n6523, A => 
                           n4567, ZN => mult_143_n4776);
   mult_143_U2396 : XNOR2_X1 port map( A => n2670, B => mult_143_n4785, ZN => 
                           SIG_in(15));
   mult_143_U2397 : AOI21_X1 port map( B1 => mult_143_n4363, B2 => n720, A => 
                           mult_143_n6526, ZN => mult_143_n4785);
   mult_143_U2412 : NOR2_X1 port map( A1 => n956, A2 => mult_143_n6536, ZN => 
                           mult_143_n4793);
   mult_143_U2413 : XNOR2_X1 port map( A => mult_143_n4795, B => mult_143_n4796
                           , ZN => SIG_in(11));
   mult_143_U2414 : AOI21_X1 port map( B1 => n4901, B2 => n4697, A => n2769, ZN
                           => mult_143_n4796);
   mult_143_U2415 : NOR2_X1 port map( A1 => n816, A2 => n2604, ZN => 
                           mult_143_n4795);
   mult_143_U2388 : NAND2_X1 port map( A1 => n4567, A2 => n953, ZN => 
                           mult_143_n4779);
   mult_143_U2389 : NOR2_X1 port map( A1 => mult_143_n6580, A2 => n727, ZN => 
                           mult_143_n4778);
   mult_143_U2368 : XNOR2_X1 port map( A => n4742, B => mult_143_n4758, ZN => 
                           SIG_in(25));
   mult_143_U2370 : NOR2_X1 port map( A1 => mult_143_n4351, A2 => 
                           mult_143_n6498, ZN => mult_143_n4758);
   mult_143_U2372 : NAND2_X1 port map( A1 => n2784, A2 => n946, ZN => 
                           mult_143_n4760);
   mult_143_U2374 : XNOR2_X1 port map( A => n1063, B => mult_143_n4762, ZN => 
                           SIG_in(23));
   mult_143_U2379 : NOR2_X1 port map( A1 => n984, A2 => mult_143_n6559, ZN => 
                           mult_143_n4762);
   mult_143_U2398 : NOR2_X1 port map( A1 => mult_143_n6526, A2 => n949, ZN => 
                           mult_143_n4786);
   mult_143_U2403 : OAI21_X1 port map( B1 => mult_143_n4791, B2 => n956, A => 
                           mult_143_n4792, ZN => mult_143_n4790);
   mult_143_U2404 : AOI21_X1 port map( B1 => n2936, B2 => n721, A => 
                           mult_143_n6536, ZN => mult_143_n4792);
   mult_143_U2392 : XNOR2_X1 port map( A => mult_143_n4781, B => n2638, ZN => 
                           SIG_in(17));
   mult_143_U2393 : AOI21_X1 port map( B1 => mult_143_n4782, B2 => n942, A => 
                           mult_143_n4339, ZN => mult_143_n4781);
   mult_143_U2394 : NOR2_X1 port map( A1 => mult_143_n4809, A2 => 
                           mult_143_n4339, ZN => mult_143_n4783);
   mult_143_U2395 : OAI21_X1 port map( B1 => mult_143_n4340, B2 => 
                           mult_143_n4784, A => mult_143_n4475, ZN => 
                           mult_143_n4782);
   mult_143_U2441 : OAI21_X1 port map( B1 => mult_143_n6496, B2 => n1698, A => 
                           n3120, ZN => mult_143_n4807);
   mult_143_U2442 : XNOR2_X1 port map( A => mult_143_n4808, B => mult_143_n6496
                           , ZN => SIG_in(2));
   mult_143_U2443 : NOR2_X1 port map( A1 => n2605, A2 => n1698, ZN => 
                           mult_143_n4808);
   mult_143_U2381 : XNOR2_X1 port map( A => n3535, B => n1699, ZN => SIG_in(21)
                           );
   mult_143_U2382 : NOR2_X1 port map( A1 => n3813, A2 => n3770, ZN => n1699);
   mult_143_U2384 : NOR2_X1 port map( A1 => mult_143_n4366, A2 => n948, ZN => 
                           mult_143_n4773);
   mult_143_U2390 : NAND2_X1 port map( A1 => mult_143_n4780, A2 => n720, ZN => 
                           mult_143_n4777);
   mult_143_U2391 : NOR2_X1 port map( A1 => mult_143_n4340, A2 => 
                           mult_143_n6518, ZN => mult_143_n4780);
   mult_143_U3733 : XNOR2_X1 port map( A => n2840, B => mult_143_n6081, ZN => 
                           mult_143_n1553);
   mult_143_U3735 : AOI21_X1 port map( B1 => n4747, B2 => n3820, A => 
                           mult_143_n6082, ZN => mult_143_n6081);
   mult_143_U3738 : AOI22_X1 port map( A1 => n4890, A2 => n3772, B1 => n4675, 
                           B2 => n2814, ZN => mult_143_n6083);
   mult_143_U2495 : AOI22_X1 port map( A1 => n3782, A2 => n3538, B1 => n3807, 
                           B2 => n3783, ZN => mult_143_n4875);
   mult_143_U3033 : NOR2_X1 port map( A1 => n3606, A2 => n3595, ZN => n1698);
   mult_143_U3111 : XNOR2_X1 port map( A => mult_143_n5558, B => mult_143_n5397
                           , ZN => n1697);
   mult_143_U3112 : XNOR2_X1 port map( A => mult_143_n5395, B => mult_143_n5396
                           , ZN => mult_143_n5558);
   mult_143_U2451 : AOI22_X1 port map( A1 => B_SIG(9), A2 => n2599, B1 => 
                           B_SIG(8), B2 => n804, ZN => mult_143_n4821);
   mult_143_U3887 : AOI222_X1 port map( A1 => n3718, A2 => n3681, B1 => n3718, 
                           B2 => n3741, C1 => n3681, C2 => n3741, ZN => n1488);
   mult_143_U3888 : XNOR2_X1 port map( A => n649, B => mult_143_n6205, ZN => 
                           mult_143_n6201);
   mult_143_U3889 : AOI21_X1 port map( B1 => B_SIG(3), B2 => n804, A => 
                           mult_143_n6206, ZN => mult_143_n6205);
   mult_143_U3890 : OAI21_X1 port map( B1 => mult_143_n4820, B2 => 
                           mult_143_n6629, A => mult_143_n6207, ZN => 
                           mult_143_n6206);
   mult_143_U3049 : AOI22_X1 port map( A1 => B_SIG(9), A2 => n772, B1 => 
                           B_SIG(8), B2 => n774, ZN => mult_143_n5491);
   mult_143_U2627 : AOI22_X1 port map( A1 => B_SIG(13), A2 => n2598, B1 => 
                           B_SIG(12), B2 => n799, ZN => mult_143_n5002);
   mult_143_U3423 : AOI21_X1 port map( B1 => n3785, B2 => n3801, A => 
                           mult_143_n5836, ZN => n1539);
   mult_143_U3424 : OAI21_X1 port map( B1 => n3666, B2 => n3659, A => 
                           mult_143_n5837, ZN => mult_143_n5836);
   mult_143_U3425 : AOI22_X1 port map( A1 => n3784, A2 => n3821, B1 => n3783, 
                           B2 => n3771, ZN => mult_143_n5837);
   mult_143_U3543 : OAI21_X1 port map( B1 => n3666, B2 => n3673, A => 
                           mult_143_n5946, ZN => mult_143_n5945);
   mult_143_U3544 : AOI22_X1 port map( A1 => n3785, A2 => n3823, B1 => n4747, 
                           B2 => n3537, ZN => mult_143_n5946);
   mult_143_U3492 : AOI21_X1 port map( B1 => n3784, B2 => n3809, A => 
                           mult_143_n5897, ZN => mult_143_n5896);
   mult_143_U3493 : OAI21_X1 port map( B1 => n3666, B2 => n3597, A => 
                           mult_143_n5898, ZN => mult_143_n5897);
   mult_143_U3494 : AOI22_X1 port map( A1 => n4695, A2 => n3808, B1 => n3783, 
                           B2 => n3536, ZN => mult_143_n5898);
   mult_143_U3897 : AOI222_X1 port map( A1 => n3740, A2 => n1065, B1 => n3740, 
                           B2 => n3719, C1 => n1065, C2 => n3719, ZN => 
                           mult_143_n1039);
   mult_143_U3898 : AOI21_X1 port map( B1 => n787, B2 => B_SIG(7), A => 
                           mult_143_n6218, ZN => mult_143_n6217);
   mult_143_U3899 : OAI21_X1 port map( B1 => mult_143_n2919, B2 => 
                           mult_143_n4828, A => mult_143_n6219, ZN => 
                           mult_143_n6218);
   mult_143_U3900 : AOI22_X1 port map( A1 => B_SIG(6), A2 => mult_143_n48, B1 
                           => B_SIG(8), B2 => n765, ZN => mult_143_n6219);
   mult_143_U3902 : XNOR2_X1 port map( A => mult_143_n6222, B => n649, ZN => 
                           n1695);
   mult_143_U3903 : AOI221_X1 port map( B1 => n2599, B2 => B_SIG(5), C1 => 
                           B_SIG(3), C2 => mult_143_n6621, A => mult_143_n6223,
                           ZN => mult_143_n6222);
   mult_143_U3904 : OAI22_X1 port map( A1 => mult_143_n3096, A2 => 
                           mult_143_n4820, B1 => n2977, B2 => n979, ZN => 
                           mult_143_n6223);
   mult_143_U3337 : OAI222_X1 port map( A1 => n2831, A2 => n2694, B1 => n2831, 
                           B2 => n2761, C1 => n2694, C2 => n2761, ZN => 
                           mult_143_n5465);
   mult_143_U2548 : AOI22_X1 port map( A1 => n3779, A2 => n3533, B1 => n3781, 
                           B2 => n3825, ZN => mult_143_n4927);
   mult_143_U3131 : XNOR2_X1 port map( A => mult_143_n5580, B => mult_143_n5581
                           , ZN => mult_143_n5216);
   mult_143_U3188 : XNOR2_X1 port map( A => mult_143_n5633, B => mult_143_n5627
                           , ZN => mult_143_n5583);
   mult_143_U3192 : XNOR2_X1 port map( A => n2884, B => mult_143_n6367, ZN => 
                           mult_143_n5633);
   mult_143_U3193 : XNOR2_X1 port map( A => mult_143_n5636, B => mult_143_n5626
                           , ZN => mult_143_n5582);
   mult_143_U3196 : XNOR2_X1 port map( A => n3047, B => mult_143_n5625, ZN => 
                           mult_143_n5636);
   mult_143_U3133 : AOI22_X1 port map( A1 => mult_143_n6388, A2 => 
                           mult_143_n5586, B1 => n730, B2 => n968, ZN => 
                           mult_143_n5585);
   mult_143_U3799 : OAI21_X1 port map( B1 => mult_143_n6098, B2 => 
                           mult_143_n6130, A => mult_143_n6118, ZN => 
                           mult_143_n6106);
   mult_143_U3800 : OAI21_X1 port map( B1 => n847, B2 => n852, A => n851, ZN =>
                           mult_143_n6118);
   mult_143_U3801 : AOI21_X1 port map( B1 => n847, B2 => n852, A => n851, ZN =>
                           mult_143_n6130);
   mult_143_U3802 : AOI21_X1 port map( B1 => mult_143_n6131, B2 => 
                           mult_143_n6002, A => mult_143_n6115, ZN => 
                           mult_143_n6098);
   mult_143_U3804 : OAI21_X1 port map( B1 => B_SIG(17), B2 => B_SIG(15), A => 
                           B_SIG(16), ZN => mult_143_n6002);
   mult_143_U3805 : OAI21_X1 port map( B1 => B_SIG(19), B2 => B_SIG(17), A => 
                           B_SIG(18), ZN => mult_143_n6131);
   mult_143_U3180 : XNOR2_X1 port map( A => n2619, B => n3816, ZN => 
                           mult_143_n5628);
   mult_143_U2523 : AOI22_X1 port map( A1 => n3784, A2 => n3807, B1 => n3783, 
                           B2 => n3538, ZN => mult_143_n4905);
   mult_143_U2553 : AOI22_X1 port map( A1 => B_SIG(9), A2 => n2598, B1 => 
                           B_SIG(8), B2 => n799, ZN => mult_143_n4933);
   mult_143_U3176 : AOI222_X1 port map( A1 => mult_143_n6367, A2 => n2884, B1 
                           => mult_143_n6367, B2 => mult_143_n5627, C1 => n2884
                           , C2 => mult_143_n5627, ZN => mult_143_n5616);
   mult_143_U3189 : NOR2_X1 port map( A1 => mult_143_n5634, A2 => 
                           mult_143_n5635, ZN => mult_143_n5627);
   mult_143_U3190 : NOR2_X1 port map( A1 => n3628, A2 => n3632, ZN => 
                           mult_143_n5635);
   mult_143_U3191 : AOI21_X1 port map( B1 => n3632, B2 => n3628, A => n3814, ZN
                           => mult_143_n5634);
   mult_143_U2994 : XNOR2_X1 port map( A => mult_143_n5417, B => mult_143_n5165
                           , ZN => n1693);
   mult_143_U2995 : AOI222_X1 port map( A1 => n714, A2 => mult_143_n6541, B1 =>
                           n714, B2 => n2615, C1 => mult_143_n6541, C2 => n2615
                           , ZN => mult_143_n5165);
   mult_143_U3671 : AOI21_X1 port map( B1 => B_SIG(19), B2 => n774, A => 
                           mult_143_n6038, ZN => mult_143_n6037);
   mult_143_U3673 : AOI22_X1 port map( A1 => B_SIG(20), A2 => n772, B1 => 
                           B_SIG(18), B2 => mult_143_n72, ZN => mult_143_n6039)
                           ;
   mult_143_U3978 : XNOR2_X1 port map( A => n1691, B => mult_143_n6279, ZN => 
                           n966);
   mult_143_U4014 : AOI221_X1 port map( B1 => B_SIG(5), B2 => n772, C1 => 
                           B_SIG(3), C2 => mult_143_n72, A => mult_143_n6304, 
                           ZN => mult_143_n6303);
   mult_143_U4015 : OAI22_X1 port map( A1 => mult_143_n3096, A2 => 
                           mult_143_n4824, B1 => n2977, B2 => n978, ZN => 
                           mult_143_n6304);
   mult_143_U3981 : AOI221_X1 port map( B1 => n804, B2 => B_SIG(7), C1 => 
                           B_SIG(6), C2 => mult_143_n6621, A => mult_143_n6283,
                           ZN => mult_143_n6282);
   mult_143_U3982 : OAI22_X1 port map( A1 => mult_143_n2919, A2 => 
                           mult_143_n4820, B1 => n886, B2 => n996, ZN => 
                           mult_143_n6283);
   mult_143_U2982 : NOR2_X1 port map( A1 => mult_143_n5206, A2 => 
                           mult_143_n5207, ZN => mult_143_n4809);
   mult_143_U3429 : AOI21_X1 port map( B1 => n2908, B2 => n3801, A => 
                           mult_143_n5842, ZN => mult_143_n5841);
   mult_143_U3744 : AOI21_X1 port map( B1 => n4890, B2 => n3820, A => 
                           mult_143_n6087, ZN => mult_143_n6086);
   mult_143_U3747 : OAI21_X1 port map( B1 => n3666, B2 => n3643, A => 
                           mult_143_n6088, ZN => mult_143_n6087);
   mult_143_U3748 : AOI22_X1 port map( A1 => n3785, A2 => n3772, B1 => n3531, 
                           B2 => n3783, ZN => mult_143_n6088);
   mult_143_U3548 : AOI21_X1 port map( B1 => n4688, B2 => n3817, A => 
                           mult_143_n5951, ZN => mult_143_n5950);
   mult_143_U3550 : AOI22_X1 port map( A1 => n3787, A2 => n3823, B1 => n4695, 
                           B2 => n3537, ZN => mult_143_n5952);
   mult_143_U3004 : NAND2_X1 port map( A1 => mult_143_n5437, A2 => n4885, ZN =>
                           mult_143_n304);
   mult_143_U3203 : NAND2_X1 port map( A1 => mult_143_n5643, A2 => 
                           mult_143_n5639, ZN => mult_143_n5170);
   mult_143_U3209 : AOI222_X1 port map( A1 => n3494, A2 => n4710, B1 => n3494, 
                           B2 => n3705, C1 => n4710, C2 => n3705, ZN => 
                           mult_143_n5643);
   mult_143_U3702 : OAI21_X1 port map( B1 => n3666, B2 => n3645, A => 
                           mult_143_n6062, ZN => mult_143_n6061);
   mult_143_U3704 : AOI22_X1 port map( A1 => n3810, A2 => n3785, B1 => n3540, 
                           B2 => n3783, ZN => mult_143_n6062);
   mult_143_U2844 : NOR2_X1 port map( A1 => n4755, A2 => n1678, ZN => 
                           mult_143_n426);
   mult_143_U3618 : XNOR2_X1 port map( A => n3796, B => n3575, ZN => n1689);
   mult_143_U3619 : AOI21_X1 port map( B1 => B_SIG(9), B2 => n774, A => 
                           mult_143_n6016, ZN => mult_143_n6015);
   mult_143_U3620 : OAI21_X1 port map( B1 => mult_143_n6627, B2 => 
                           mult_143_n4824, A => mult_143_n6017, ZN => 
                           mult_143_n6016);
   mult_143_U3621 : AOI22_X1 port map( A1 => B_SIG(10), A2 => n772, B1 => 
                           B_SIG(8), B2 => mult_143_n72, ZN => mult_143_n6017);
   mult_143_U3407 : AOI21_X1 port map( B1 => B_SIG(13), B2 => mult_143_n2, A =>
                           mult_143_n5821, ZN => mult_143_n5820);
   mult_143_U3408 : OAI21_X1 port map( B1 => mult_143_n5124, B2 => 
                           mult_143_n3010, A => mult_143_n5822, ZN => 
                           mult_143_n5821);
   mult_143_U3410 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n1030, B1 => 
                           B_SIG(12), B2 => mult_143_n3245, ZN => 
                           mult_143_n5822);
   mult_143_U3588 : AOI21_X1 port map( B1 => n3827, B2 => n4664, A => 
                           mult_143_n5988, ZN => mult_143_n5987);
   mult_143_U3589 : OAI21_X1 port map( B1 => n3594, B2 => n3665, A => 
                           mult_143_n5989, ZN => mult_143_n5988);
   mult_143_U3590 : AOI22_X1 port map( A1 => n3800, A2 => n4656, B1 => n3767, 
                           B2 => n4845, ZN => mult_143_n5989);
   mult_143_U3025 : NOR2_X1 port map( A1 => mult_143_n5436, A2 => 
                           mult_143_n5437, ZN => n948);
   mult_143_U3027 : XNOR2_X1 port map( A => n4839, B => mult_143_n5463, ZN => 
                           mult_143_n5461);
   mult_143_U3031 : AOI222_X1 port map( A1 => n1648, A2 => n3555, B1 => n3555, 
                           B2 => n3737, C1 => n1648, C2 => n3737, ZN => 
                           mult_143_n5436);
   mult_143_U3306 : XNOR2_X1 port map( A => mult_143_n5740, B => mult_143_n5741
                           , ZN => n1688);
   mult_143_U3477 : AOI21_X1 port map( B1 => B_SIG(12), B2 => n1031, A => 
                           mult_143_n5882, ZN => mult_143_n5881);
   mult_143_U3478 : OAI21_X1 port map( B1 => mult_143_n5859, B2 => 
                           mult_143_n3010, A => mult_143_n5883, ZN => 
                           mult_143_n5882);
   mult_143_U3530 : AOI21_X1 port map( B1 => n3817, B2 => n4845, A => 
                           mult_143_n5933, ZN => mult_143_n5932);
   mult_143_U3531 : OAI21_X1 port map( B1 => n3673, B2 => n3665, A => 
                           mult_143_n5934, ZN => mult_143_n5933);
   mult_143_U2930 : XNOR2_X1 port map( A => n2618, B => n2766, ZN => 
                           mult_143_n5351);
   mult_143_U2825 : NAND2_X1 port map( A1 => mult_143_n5206, A2 => 
                           mult_143_n5207, ZN => mult_143_n344);
   mult_143_U3265 : XNOR2_X1 port map( A => n3736, B => n3523, ZN => n1687);
   mult_143_U3266 : XNOR2_X1 port map( A => mult_143_n5700, B => mult_143_n5701
                           , ZN => mult_143_n5698);
   mult_143_U3286 : XNOR2_X1 port map( A => mult_143_n5716, B => mult_143_n6555
                           , ZN => mult_143_n5700);
   mult_143_U3287 : XNOR2_X1 port map( A => n2717, B => mult_143_n6554, ZN => 
                           mult_143_n5716);
   mult_143_U3275 : XNOR2_X1 port map( A => mult_143_n5707, B => mult_143_n5706
                           , ZN => n1686);
   mult_143_U3276 : AOI21_X1 port map( B1 => mult_143_n5708, B2 => 
                           mult_143_n5709, A => mult_143_n5710, ZN => 
                           mult_143_n5706);
   mult_143_U3277 : NOR2_X1 port map( A1 => mult_143_n5709, A2 => 
                           mult_143_n5708, ZN => mult_143_n5710);
   mult_143_U3317 : AOI222_X1 port map( A1 => n717, A2 => n4838, B1 => n717, B2
                           => n2721, C1 => n4838, C2 => n2721, ZN => 
                           mult_143_n5470);
   mult_143_U3318 : AOI222_X1 port map( A1 => n2665, A2 => n3058, B1 => n2665, 
                           B2 => n3803, C1 => n3058, C2 => n3803, ZN => 
                           mult_143_n5747);
   mult_143_U3195 : AOI21_X1 port map( B1 => mult_143_n5228, B2 => n2767, A => 
                           n2668, ZN => mult_143_n5637);
   mult_143_U3854 : OAI21_X1 port map( B1 => mult_143_n4828, B2 => 
                           mult_143_n6629, A => mult_143_n6172, ZN => 
                           mult_143_n6171);
   mult_143_U3849 : AOI21_X1 port map( B1 => B_SIG(5), B2 => mult_143_n36, A =>
                           mult_143_n6166, ZN => mult_143_n6165);
   mult_143_U3850 : OAI21_X1 port map( B1 => mult_143_n2798, B2 => 
                           mult_143_n4848, A => mult_143_n6167, ZN => 
                           mult_143_n6166);
   mult_143_U3851 : AOI22_X1 port map( A1 => B_SIG(7), A2 => n755, B1 => 
                           B_SIG(6), B2 => n1023, ZN => mult_143_n6167);
   mult_143_U2586 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n2598, B1 => 
                           B_SIG(9), B2 => mult_143_n96, ZN => mult_143_n4961);
   mult_143_U3245 : XNOR2_X1 port map( A => mult_143_n5682, B => n3734, ZN => 
                           mult_143_n5188);
   mult_143_U3246 : XNOR2_X1 port map( A => mult_143_n5684, B => mult_143_n5683
                           , ZN => n1685);
   mult_143_U3285 : AOI222_X1 port map( A1 => mult_143_n2759, A2 => 
                           mult_143_n6367, B1 => mult_143_n2759, B2 => 
                           mult_143_n6368, C1 => mult_143_n6367, C2 => 
                           mult_143_n6368, ZN => mult_143_n5685);
   mult_143_U3247 : XNOR2_X1 port map( A => n1471, B => n3733, ZN => 
                           mult_143_n5682);
   mult_143_U3248 : XNOR2_X1 port map( A => mult_143_n5688, B => mult_143_n5687
                           , ZN => n1684);
   mult_143_U3249 : XNOR2_X1 port map( A => mult_143_n5689, B => mult_143_n5690
                           , ZN => mult_143_n5687);
   mult_143_U3271 : XNOR2_X1 port map( A => mult_143_n5703, B => mult_143_n6563
                           , ZN => mult_143_n5690);
   mult_143_U3272 : XNOR2_X1 port map( A => mult_143_n6367, B => n2719, ZN => 
                           mult_143_n5703);
   mult_143_U3273 : XNOR2_X1 port map( A => mult_143_n5704, B => mult_143_n5705
                           , ZN => mult_143_n5689);
   mult_143_U3274 : XNOR2_X1 port map( A => n2869, B => n4878, ZN => 
                           mult_143_n5704);
   mult_143_U3258 : XNOR2_X1 port map( A => mult_143_n6368, B => mult_143_n5692
                           , ZN => mult_143_n5679);
   mult_143_U2641 : AOI222_X1 port map( A1 => n1629, A2 => n3099, B1 => n1629, 
                           B2 => n666, C1 => n3099, C2 => n666, ZN => 
                           mult_143_n759);
   mult_143_U3878 : AOI21_X1 port map( B1 => mult_143_n3228, B2 => B_SIG(10), A
                           => mult_143_n6196, ZN => mult_143_n6195);
   mult_143_U3879 : OAI21_X1 port map( B1 => mult_143_n6626, B2 => 
                           mult_143_n5859, A => mult_143_n6197, ZN => 
                           mult_143_n6196);
   mult_143_U3880 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n1031, B1 => 
                           B_SIG(12), B2 => n1026, ZN => mult_143_n6197);
   mult_143_U3211 : XNOR2_X1 port map( A => mult_143_n5660, B => mult_143_n5661
                           , ZN => mult_143_n5654);
   mult_143_U3212 : AOI22_X1 port map( A1 => mult_143_n6369, A2 => n3590, B1 =>
                           n4593, B2 => n969, ZN => mult_143_n5661);
   mult_143_U3213 : XNOR2_X1 port map( A => mult_143_n5662, B => mult_143_n5663
                           , ZN => mult_143_n5653);
   mult_143_U3214 : AOI22_X1 port map( A1 => mult_143_n6543, A2 => n994, B1 => 
                           n4690, B2 => n970, ZN => mult_143_n5663);
   mult_143_U3146 : XNOR2_X1 port map( A => mult_143_n6610, B => mult_143_n5601
                           , ZN => mult_143_n5600);
   mult_143_U3591 : AOI21_X1 port map( B1 => n4736, B2 => n4665, A => 
                           mult_143_n5991, ZN => n1538);
   mult_143_U3593 : AOI22_X1 port map( A1 => n3800, A2 => n4664, B1 => n3782, 
                           B2 => n4656, ZN => mult_143_n5992);
   mult_143_U3639 : XNOR2_X1 port map( A => n4760, B => mult_143_n6023, ZN => 
                           n1040);
   mult_143_U3644 : AOI21_X1 port map( B1 => n4736, B2 => n3819, A => 
                           mult_143_n6024, ZN => mult_143_n6023);
   mult_143_U3646 : AOI22_X1 port map( A1 => n3766, A2 => n3533, B1 => n4675, 
                           B2 => n3825, ZN => mult_143_n6025);
   mult_143_U2887 : AOI222_X1 port map( A1 => n3617, A2 => n3623, B1 => n3617, 
                           B2 => n3639, C1 => n3623, C2 => n3639, ZN => 
                           mult_143_n5294);
   mult_143_U2488 : AOI22_X1 port map( A1 => n3779, A2 => n3538, B1 => n3781, 
                           B2 => n4848, ZN => mult_143_n4864);
   mult_143_U3416 : AOI22_X1 port map( A1 => n3800, A2 => n3771, B1 => n4736, 
                           B2 => n3762, ZN => mult_143_n5828);
   mult_143_U3442 : NOR3_X1 port map( A1 => A_SIG(0), A2 => A_SIG(1), A3 => 
                           n536, ZN => mult_143_n3239);
   mult_143_U3449 : AOI22_X1 port map( A1 => A_SIG(2), A2 => A_SIG(1), B1 => 
                           n639, B2 => n536, ZN => mult_143_n5853);
   mult_143_U3575 : AOI22_X1 port map( A1 => n3800, A2 => n3798, B1 => n3781, 
                           B2 => n3807, ZN => mult_143_n5976);
   mult_143_U3627 : AOI21_X1 port map( B1 => B_SIG(12), B2 => n774, A => 
                           mult_143_n6019, ZN => mult_143_n6018);
   mult_143_U3637 : OAI21_X1 port map( B1 => mult_143_n4824, B2 => 
                           mult_143_n3010, A => mult_143_n6020, ZN => 
                           mult_143_n6019);
   mult_143_U2794 : AOI222_X1 port map( A1 => n3605, A2 => n3730, B1 => n3605, 
                           B2 => n3509, C1 => n3730, C2 => n3509, ZN => 
                           mult_143_n5168);
   mult_143_U2795 : AOI222_X1 port map( A1 => mult_143_n5160, A2 => 
                           mult_143_n5161, B1 => mult_143_n5160, B2 => 
                           mult_143_n5159, C1 => mult_143_n5159, C2 => 
                           mult_143_n5161, ZN => n1486);
   mult_143_U2796 : XNOR2_X1 port map( A => mult_143_n5174, B => mult_143_n5175
                           , ZN => mult_143_n5159);
   mult_143_U2797 : AOI22_X1 port map( A1 => mult_143_n6564, A2 => n991, B1 => 
                           n4949, B2 => mult_143_n4355, ZN => mult_143_n5175);
   mult_143_U2798 : XNOR2_X1 port map( A => n3059, B => mult_143_n5176, ZN => 
                           mult_143_n5161);
   mult_143_U2799 : AOI22_X1 port map( A1 => mult_143_n6374, A2 => n3099, B1 =>
                           n2864, B2 => n957, ZN => mult_143_n5176);
   mult_143_U2989 : XNOR2_X1 port map( A => n2600, B => mult_143_n6473, ZN => 
                           mult_143_n5178);
   mult_143_U2991 : XNOR2_X1 port map( A => mult_143_n5416, B => n2691, ZN => 
                           mult_143_n5177);
   mult_143_U2992 : XNOR2_X1 port map( A => n2727, B => n2669, ZN => 
                           mult_143_n5416);
   mult_143_U2801 : XNOR2_X1 port map( A => mult_143_n5180, B => mult_143_n5179
                           , ZN => n1681);
   mult_143_U2802 : XNOR2_X1 port map( A => mult_143_n5181, B => mult_143_n5182
                           , ZN => mult_143_n5179);
   mult_143_U3219 : XNOR2_X1 port map( A => n2634, B => n2778, ZN => 
                           mult_143_n5664);
   mult_143_U3220 : AOI21_X1 port map( B1 => n957, B2 => n2864, A => 
                           mult_143_n5665, ZN => mult_143_n5181);
   mult_143_U3221 : AOI21_X1 port map( B1 => mult_143_n6374, B2 => n3099, A => 
                           n3059, ZN => mult_143_n5665);
   mult_143_U3229 : XNOR2_X1 port map( A => mult_143_n5667, B => mult_143_n5668
                           , ZN => mult_143_n5186);
   mult_143_U3230 : AOI22_X1 port map( A1 => mult_143_n6598, A2 => n3678, B1 =>
                           n4616, B2 => n971, ZN => mult_143_n5668);
   mult_143_U3540 : AOI22_X1 port map( A1 => n3800, A2 => n3537, B1 => n3782, 
                           B2 => n3823, ZN => mult_143_n5943);
   mult_143_U3483 : AOI21_X1 port map( B1 => n4736, B2 => n3809, A => 
                           mult_143_n5888, ZN => mult_143_n5887);
   mult_143_U3485 : AOI22_X1 port map( A1 => n3800, A2 => n3536, B1 => n3782, 
                           B2 => n3808, ZN => mult_143_n5889);
   mult_143_U2505 : AOI222_X1 port map( A1 => n1623, A2 => n3691, B1 => n1623, 
                           B2 => n1621, C1 => n1621, C2 => n3691, ZN => 
                           mult_143_n901);
   mult_143_U2512 : AOI21_X1 port map( B1 => mult_143_n72, B2 => B_SIG(10), A 
                           => mult_143_n4894, ZN => mult_143_n4893);
   mult_143_U2513 : OAI21_X1 port map( B1 => mult_143_n6626, B2 => 
                           mult_143_n4824, A => mult_143_n4895, ZN => 
                           mult_143_n4894);
   mult_143_U2514 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n774, B1 => 
                           B_SIG(12), B2 => n772, ZN => mult_143_n4895);
   mult_143_U3918 : AOI222_X1 port map( A1 => n1670, A2 => n3729, B1 => n1670, 
                           B2 => n1669, C1 => n3729, C2 => n1669, ZN => 
                           mult_143_n1027);
   mult_143_U3937 : XNOR2_X1 port map( A => n649, B => mult_143_n6246, ZN => 
                           n1679);
   mult_143_U3938 : AOI21_X1 port map( B1 => B_SIG(5), B2 => n804, A => 
                           mult_143_n6247, ZN => mult_143_n6246);
   mult_143_U3939 : OAI21_X1 port map( B1 => mult_143_n4820, B2 => 
                           mult_143_n2800, A => mult_143_n6248, ZN => 
                           mult_143_n6247);
   mult_143_U3942 : AOI21_X1 port map( B1 => B_SIG(10), B2 => mult_143_n36, A 
                           => mult_143_n6251, ZN => mult_143_n6250);
   mult_143_U3943 : OAI21_X1 port map( B1 => mult_143_n6626, B2 => 
                           mult_143_n4848, A => mult_143_n6252, ZN => 
                           mult_143_n6251);
   mult_143_U3944 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n1023, B1 => 
                           B_SIG(12), B2 => n755, ZN => mult_143_n6252);
   mult_143_U2923 : NOR2_X1 port map( A1 => mult_143_n5343, A2 => 
                           mult_143_n5344, ZN => mult_143_n5333);
   mult_143_U2924 : NOR2_X1 port map( A1 => n3635, A2 => n3637, ZN => 
                           mult_143_n5344);
   mult_143_U2925 : AOI21_X1 port map( B1 => n3637, B2 => n3635, A => n1758, ZN
                           => mult_143_n5343);
   mult_143_U3120 : AOI222_X1 port map( A1 => n967, A2 => n992, B1 => n967, B2 
                           => mult_143_n5552, C1 => n992, C2 => mult_143_n5552,
                           ZN => mult_143_n5559);
   mult_143_U3138 : XNOR2_X1 port map( A => mult_143_n5589, B => n3619, ZN => 
                           mult_143_n5564);
   mult_143_U3139 : XNOR2_X1 port map( A => n3630, B => n4633, ZN => 
                           mult_143_n5589);
   mult_143_U3140 : NOR2_X1 port map( A1 => mult_143_n5590, A2 => 
                           mult_143_n5591, ZN => mult_143_n5562);
   mult_143_U3142 : AOI21_X1 port map( B1 => n3107, B2 => mult_143_n6408, A => 
                           n2608, ZN => mult_143_n5590);
   mult_143_U3124 : XNOR2_X1 port map( A => mult_143_n5572, B => mult_143_n5571
                           , ZN => mult_143_n5569);
   mult_143_U3143 : XNOR2_X1 port map( A => mult_143_n5592, B => mult_143_n6401
                           , ZN => mult_143_n5572);
   mult_143_U3184 : XNOR2_X1 port map( A => mult_143_n6611, B => n1606, ZN => 
                           mult_143_n5594);
   mult_143_U3109 : XNOR2_X1 port map( A => mult_143_n5552, B => mult_143_n5553
                           , ZN => mult_143_n5481);
   mult_143_U3110 : AOI22_X1 port map( A1 => mult_143_n6406, A2 => n992, B1 => 
                           mult_143_n6407, B2 => n967, ZN => mult_143_n5553);
   mult_143_U3121 : XNOR2_X1 port map( A => n3629, B => mult_143_n5567, ZN => 
                           mult_143_n5552);
   mult_143_U3105 : XNOR2_X1 port map( A => n2622, B => mult_143_n5550, ZN => 
                           mult_143_n5478);
   mult_143_U3952 : OAI21_X1 port map( B1 => mult_143_n6080, B2 => 
                           mult_143_n6258, A => mult_143_n6259, ZN => 
                           mult_143_n6127);
   mult_143_U3954 : AOI21_X1 port map( B1 => n891, B2 => n882, A => n886, ZN =>
                           mult_143_n6080);
   mult_143_U2640 : AOI22_X1 port map( A1 => n3792, A2 => mult_143_n1532, B1 =>
                           n666, B2 => n3768, ZN => mult_143_n5015);
   mult_143_U2643 : OAI21_X1 port map( B1 => n3643, B2 => n3667, A => 
                           mult_143_n5018, ZN => mult_143_n5017);
   mult_143_U2846 : NAND2_X1 port map( A1 => mult_143_n5243, A2 => n1615, ZN =>
                           mult_143_n5242);
   mult_143_U2847 : NAND2_X1 port map( A1 => mult_143_n5239, A2 => n4573, ZN =>
                           mult_143_n5243);
   mult_143_U2951 : NAND2_X1 port map( A1 => n3609, A2 => n3507, ZN => 
                           mult_143_n5239);
   mult_143_U2952 : AOI222_X1 port map( A1 => n702, A2 => mult_143_n5251, B1 =>
                           n702, B2 => mult_143_n5252, C1 => mult_143_n5252, C2
                           => mult_143_n5251, ZN => n1483);
   mult_143_U2953 : XNOR2_X1 port map( A => mult_143_n5379, B => mult_143_n5380
                           , ZN => mult_143_n5252);
   mult_143_U2954 : XNOR2_X1 port map( A => mult_143_n5382, B => n2705, ZN => 
                           mult_143_n5251);
   mult_143_U2955 : XNOR2_X1 port map( A => mult_143_n6427, B => n2877, ZN => 
                           mult_143_n5382);
   mult_143_U2956 : OAI222_X1 port map( A1 => n4781, A2 => n2618, B1 => n4781, 
                           B2 => n2766, C1 => n2766, C2 => n2618, ZN => 
                           mult_143_n5250);
   mult_143_U2959 : XNOR2_X1 port map( A => mult_143_n6573, B => mult_143_n5384
                           , ZN => mult_143_n5380);
   mult_143_U2960 : AOI22_X1 port map( A1 => n2695, A2 => mult_143_n6572, B1 =>
                           n986, B2 => n1657, ZN => mult_143_n5384);
   mult_143_U2963 : XNOR2_X1 port map( A => mult_143_n5385, B => n3093, ZN => 
                           mult_143_n5377);
   mult_143_U2964 : XNOR2_X1 port map( A => mult_143_n6421, B => n2711, ZN => 
                           mult_143_n5385);
   mult_143_U2965 : XNOR2_X1 port map( A => mult_143_n5387, B => n2888, ZN => 
                           mult_143_n5376);
   mult_143_U3050 : XNOR2_X1 port map( A => mult_143_n5492, B => n3773, ZN => 
                           n1677);
   mult_143_U3052 : OAI21_X1 port map( B1 => n3664, B2 => n3594, A => 
                           mult_143_n5494, ZN => mult_143_n5493);
   mult_143_U3053 : AOI22_X1 port map( A1 => n3827, A2 => n3767, B1 => n4845, 
                           B2 => n4656, ZN => mult_143_n5494);
   mult_143_U3345 : NOR2_X1 port map( A1 => mult_143_n5770, A2 => 
                           mult_143_n5771, ZN => mult_143_n5463);
   mult_143_U3346 : NOR2_X1 port map( A1 => mult_143_n4490, A2 => n3824, ZN => 
                           mult_143_n5771);
   mult_143_U3347 : AOI21_X1 port map( B1 => n3824, B2 => mult_143_n4490, A => 
                           mult_143_n706, ZN => mult_143_n5770);
   mult_143_U3348 : XNOR2_X1 port map( A => mult_143_n5772, B => mult_143_n4490
                           , ZN => mult_143_n5462);
   mult_143_U3349 : XNOR2_X1 port map( A => n2696, B => n3065, ZN => 
                           mult_143_n5772);
   mult_143_U3321 : AOI222_X1 port map( A1 => n2624, A2 => n4754, B1 => n2624, 
                           B2 => n2666, C1 => n2666, C2 => n4754, ZN => 
                           mult_143_n5728);
   mult_143_U3156 : XNOR2_X1 port map( A => mult_143_n6381, B => mult_143_n5609
                           , ZN => n1676);
   mult_143_U3158 : XNOR2_X1 port map( A => mult_143_n6382, B => n3116, ZN => 
                           mult_143_n5611);
   mult_143_U3159 : AOI222_X1 port map( A1 => n4744, A2 => n2759, B1 => n4744, 
                           B2 => mult_143_n5613, C1 => n2759, C2 => 
                           mult_143_n5613, ZN => n1482);
   mult_143_U3171 : XNOR2_X1 port map( A => mult_143_n5623, B => n2737, ZN => 
                           mult_143_n5613);
   mult_143_U3161 : AOI222_X1 port map( A1 => mult_143_n6385, A2 => n3062, B1 
                           => mult_143_n6385, B2 => n2737, C1 => n3062, C2 => 
                           n2737, ZN => mult_143_n5424);
   mult_143_U3163 : AOI222_X1 port map( A1 => n2619, A2 => n3816, B1 => n3816, 
                           B2 => mult_143_n5619, C1 => n2619, C2 => 
                           mult_143_n5619, ZN => mult_143_n5418);
   mult_143_U3177 : NOR2_X1 port map( A1 => mult_143_n5629, A2 => 
                           mult_143_n5630, ZN => mult_143_n5619);
   mult_143_U3178 : NOR2_X1 port map( A1 => n3815, A2 => n3627, ZN => 
                           mult_143_n5630);
   mult_143_U3179 : AOI21_X1 port map( B1 => n3627, B2 => n3815, A => n3631, ZN
                           => mult_143_n5629);
   mult_143_U2510 : OAI21_X1 port map( B1 => mult_143_n4891, B2 => 
                           mult_143_n2800, A => mult_143_n4892, ZN => 
                           mult_143_n4890);
   mult_143_U2447 : AOI222_X1 port map( A1 => n1617, A2 => n3689, B1 => n1617, 
                           B2 => n3651, C1 => n3689, C2 => n3651, ZN => n967);
   mult_143_U2452 : AOI21_X1 port map( B1 => n774, B2 => B_SIG(5), A => 
                           mult_143_n4823, ZN => mult_143_n4822);
   mult_143_U2453 : OAI21_X1 port map( B1 => mult_143_n4824, B2 => 
                           mult_143_n2800, A => mult_143_n4825, ZN => 
                           mult_143_n4823);
   mult_143_U2455 : AOI21_X1 port map( B1 => mult_143_n48, B2 => B_SIG(10), A 
                           => mult_143_n4827, ZN => mult_143_n4826);
   mult_143_U2456 : OAI21_X1 port map( B1 => mult_143_n6626, B2 => 
                           mult_143_n4828, A => mult_143_n4829, ZN => 
                           mult_143_n4827);
   mult_143_U2457 : AOI22_X1 port map( A1 => B_SIG(11), A2 => n787, B1 => 
                           B_SIG(12), B2 => n765, ZN => mult_143_n4829);
   mult_143_U2902 : NOR2_X1 port map( A1 => mult_143_n5327, A2 => 
                           mult_143_n5328, ZN => mult_143_n5320);
   mult_143_U2903 : NOR2_X1 port map( A1 => n1751, A2 => n1739, ZN => 
                           mult_143_n5328);
   mult_143_U2904 : AOI21_X1 port map( B1 => n1739, B2 => n1751, A => n1740, ZN
                           => mult_143_n5327);
   mult_143_U3907 : AOI221_X1 port map( B1 => B_SIG(3), B2 => n772, C1 => 
                           B_SIG(1), C2 => mult_143_n72, A => mult_143_n6229, 
                           ZN => mult_143_n6228);
   mult_143_U3909 : OAI22_X1 port map( A1 => mult_143_n6630, A2 => 
                           mult_143_n4824, B1 => n910, B2 => n978, ZN => 
                           mult_143_n6229);
   mult_143_U3916 : OAI22_X1 port map( A1 => n910, A2 => n977, B1 => 
                           mult_143_n4824, B2 => n2817, ZN => mult_143_n6234);
   mult_143_U3961 : XNOR2_X1 port map( A => n3520, B => n1671, ZN => n962);
   mult_143_U3967 : XNOR2_X1 port map( A => n649, B => mult_143_n6267, ZN => 
                           mult_143_n6264);
   mult_143_U3968 : AOI21_X1 port map( B1 => B_SIG(5), B2 => mult_143_n6621, A 
                           => mult_143_n6268, ZN => mult_143_n6267);
   mult_143_U3969 : OAI21_X1 port map( B1 => mult_143_n2798, B2 => 
                           mult_143_n4820, A => mult_143_n6269, ZN => 
                           mult_143_n6268);
   mult_143_U3970 : AOI22_X1 port map( A1 => B_SIG(7), A2 => n2599, B1 => 
                           B_SIG(6), B2 => n804, ZN => mult_143_n6269);
   mult_143_U3973 : OAI21_X1 port map( B1 => mult_143_n4824, B2 => 
                           mult_143_n6629, A => mult_143_n6275, ZN => 
                           mult_143_n6274);
   mult_143_U2889 : OAI222_X1 port map( A1 => mult_143_n5315, A2 => n3615, B1 
                           => mult_143_n5315, B2 => n2703, C1 => n3615, C2 => 
                           n2703, ZN => mult_143_n5316);
   mult_143_U3872 : AOI21_X1 port map( B1 => n787, B2 => B_SIG(5), A => 
                           mult_143_n6190, ZN => mult_143_n6189);
   mult_143_U3873 : OAI21_X1 port map( B1 => mult_143_n4828, B2 => 
                           mult_143_n2800, A => mult_143_n6191, ZN => 
                           mult_143_n6190);
   mult_143_U2525 : AOI22_X1 port map( A1 => n3567, A2 => n3724, B1 => n4599, 
                           B2 => n4604, ZN => mult_143_n886);
   mult_143_U2527 : XNOR2_X1 port map( A => n748, B => mult_143_n4908, ZN => 
                           n1674);
   mult_143_U2528 : AOI21_X1 port map( B1 => B_SIG(5), B2 => mult_143_n96, A =>
                           mult_143_n4909, ZN => mult_143_n4908);
   mult_143_U2529 : OAI21_X1 port map( B1 => mult_143_n2798, B2 => 
                           mult_143_n4891, A => mult_143_n4910, ZN => 
                           mult_143_n4909);
   mult_143_U2530 : AOI22_X1 port map( A1 => B_SIG(7), A2 => n2598, B1 => 
                           B_SIG(6), B2 => n799, ZN => mult_143_n4910);
   mult_143_U3584 : OAI21_X1 port map( B1 => mult_143_n6629, B2 => 
                           mult_143_n4467, A => mult_143_n1910, ZN => n1535);
   mult_143_U3975 : XNOR2_X1 port map( A => n631, B => mult_143_n6276, ZN => 
                           mult_143_n6629);
   mult_143_U3976 : OAI21_X1 port map( B1 => B_SIG(3), B2 => B_SIG(4), A => 
                           mult_143_n6277, ZN => mult_143_n6276);
   mult_143_U3977 : NAND2_X1 port map( A1 => B_SIG(3), A2 => B_SIG(4), ZN => 
                           mult_143_n6277);
   mult_143_U2550 : AOI222_X1 port map( A1 => n1627, A2 => n1626, B1 => n1627, 
                           B2 => n3826, C1 => n1626, C2 => n3826, ZN => n971);
   mult_143_U2532 : AOI22_X1 port map( A1 => n3566, A2 => n1673, B1 => n2718, 
                           B2 => n4605, ZN => n961);
   mult_143_U2534 : XNOR2_X1 port map( A => n2840, B => n3521, ZN => n1673);
   mult_143_U2535 : AOI221_X1 port map( B1 => n799, B2 => B_SIG(7), C1 => 
                           B_SIG(6), C2 => mult_143_n96, A => mult_143_n4914, 
                           ZN => mult_143_n4913);
   mult_143_U2536 : OAI22_X1 port map( A1 => mult_143_n2919, A2 => 
                           mult_143_n4891, B1 => n886, B2 => n997, ZN => 
                           mult_143_n4914);
   mult_143_U3991 : AOI21_X1 port map( B1 => B_SIG(8), B2 => B_SIG(7), A => 
                           mult_143_n6291, ZN => mult_143_n6285);
   mult_143_U3992 : NOR2_X1 port map( A1 => B_SIG(7), A2 => B_SIG(8), ZN => 
                           mult_143_n6291);
   mult_143_U4389 : OAI21_X1 port map( B1 => n1068, B2 => mult_143_n4467, A => 
                           mult_143_n1909, ZN => n1534);
   mult_143_U4207 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(5), B1 => 
                           mult_143_n4468, B2 => B_SIG(4), C1 => mult_143_n4468
                           , C2 => B_SIG(3), ZN => mult_143_n1909);
   mult_143_U3836 : OAI21_X1 port map( B1 => mult_143_n6630, B2 => 
                           mult_143_n4828, A => mult_143_n6156, ZN => 
                           mult_143_n6155);
   mult_143_U3837 : AOI22_X1 port map( A1 => B_SIG(1), A2 => mult_143_n48, B1 
                           => B_SIG(2), B2 => n787, ZN => mult_143_n6156);
   mult_143_U3021 : NAND2_X1 port map( A1 => mult_143_n5446, A2 => 
                           mult_143_n5445, ZN => mult_143_n3075);
   mult_143_U4056 : OAI21_X1 port map( B1 => mult_143_n2800, B2 => 
                           mult_143_n4467, A => mult_143_n1908, ZN => 
                           mult_143_n1537);
   mult_143_U4252 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(6), B1 => 
                           mult_143_n4468, B2 => B_SIG(5), C1 => mult_143_n4468
                           , C2 => B_SIG(4), ZN => mult_143_n1908);
   mult_143_U3941 : AOI22_X1 port map( A1 => B_SIG(5), A2 => n895, B1 => 
                           B_SIG(6), B2 => n2978, ZN => mult_143_n6249);
   mult_143_U2554 : AOI21_X1 port map( B1 => B_SIG(11), B2 => n1027, A => 
                           mult_143_n4935, ZN => mult_143_n4934);
   mult_143_U2555 : OAI21_X1 port map( B1 => mult_143_n6626, B2 => 
                           mult_143_n4842, A => mult_143_n4936, ZN => 
                           mult_143_n4935);
   mult_143_U2556 : AOI22_X1 port map( A1 => mult_143_n74, A2 => B_SIG(12), B1 
                           => mult_143_n84, B2 => B_SIG(10), ZN => 
                           mult_143_n4936);
   mult_143_U3949 : OAI21_X1 port map( B1 => B_SIG(11), B2 => B_SIG(12), A => 
                           mult_143_n6257, ZN => mult_143_n6256);
   mult_143_U3950 : NAND2_X1 port map( A1 => B_SIG(11), A2 => B_SIG(12), ZN => 
                           mult_143_n6257);
   mult_143_U3656 : AOI222_X1 port map( A1 => mult_143_n4156, A2 => B_SIG(4), 
                           B1 => mult_143_n4275, B2 => B_SIG(3), C1 => 
                           mult_143_n4217, C2 => B_SIG(2), ZN => mult_143_n1863
                           );
   mult_143_U4212 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(4), B1 => 
                           mult_143_n4468, B2 => B_SIG(3), C1 => mult_143_n4468
                           , C2 => B_SIG(2), ZN => mult_143_n1910);
   mult_143_U3664 : AOI222_X1 port map( A1 => mult_143_n4154, A2 => B_SIG(14), 
                           B1 => mult_143_n4273, B2 => B_SIG(13), C1 => 
                           mult_143_n4215, C2 => B_SIG(12), ZN => 
                           mult_143_n1853);
   mult_143_U3908 : OAI21_X1 port map( B1 => n2817, B2 => mult_143_n4467, A => 
                           mult_143_n1912, ZN => mult_143_n922);
   mult_143_U4275 : OAI21_X1 port map( B1 => mult_143_n4467, B2 => n629, A => 
                           mult_143_n2743, ZN => n1533);
   mult_143_U2595 : AOI222_X1 port map( A1 => mult_143_n1536, A2 => n693, B1 =>
                           mult_143_n1536, B2 => n686, C1 => n693, C2 => n686, 
                           ZN => n1481);
   mult_143_U3825 : OAI21_X1 port map( B1 => mult_143_n4467, B2 => 
                           mult_143_n2458, A => mult_143_n1127, ZN => 
                           mult_143_n938);
   mult_143_U3647 : AOI22_X1 port map( A1 => mult_143_n4319, A2 => B_SIG(1), B1
                           => mult_143_n4201, B2 => B_SIG(0), ZN => 
                           mult_143_n1123);
   mult_143_U3409 : AOI22_X1 port map( A1 => mult_143_n4468, A2 => B_SIG(0), B1
                           => n748, B2 => B_SIG(1), ZN => mult_143_n1127);
   mult_143_U3711 : AOI222_X1 port map( A1 => n748, A2 => B_SIG(2), B1 => 
                           mult_143_n4468, B2 => B_SIG(1), C1 => mult_143_n4468
                           , C2 => B_SIG(0), ZN => mult_143_n1912);
   mult_143_U4674 : OAI33_X1 port map( A1 => B_SIG(3), A2 => n2823, A3 => n2977
                           , B1 => n909, B2 => n631, B3 => B_SIG(4), ZN => 
                           mult_143_n6307);
   mult_143_U4672 : XOR2_X1 port map( A => A_SIG(17), B => mult_143_n6303, Z =>
                           n1672);
   mult_143_U4670 : XOR2_X1 port map( A => A_SIG(20), B => mult_143_n6297, Z =>
                           mult_143_n4844);
   mult_143_U4669 : XOR2_X1 port map( A => mult_143_n6294, B => A_SIG(20), Z =>
                           mult_143_n6265);
   mult_143_U4667 : NAND3_X1 port map( A1 => B_SIG(5), A2 => B_SIG(7), A3 => 
                           mult_143_n6272, ZN => mult_143_n6287);
   mult_143_U4665 : XOR2_X1 port map( A => n3723, B => n3682, Z => 
                           mult_143_n6279);
   mult_143_U4664 : XOR2_X1 port map( A => A_SIG(17), B => mult_143_n6273, Z =>
                           mult_143_n6263);
   mult_143_U4661 : XOR2_X1 port map( A => n3722, B => n3725, Z => n1671);
   mult_143_U4658 : XOR2_X1 port map( A => n3569, B => n3793, Z => n1670);
   mult_143_U4651 : XOR2_X1 port map( A => A_SIG(17), B => mult_143_n6233, Z =>
                           n1668);
   mult_143_U4649 : XOR2_X1 port map( A => A_SIG(17), B => mult_143_n6228, Z =>
                           n1667);
   mult_143_U4647 : XOR2_X1 port map( A => mult_143_n6217, B => A_SIG(11), Z =>
                           n1666);
   mult_143_U4645 : XOR2_X1 port map( A => mult_143_n6210, B => A_SIG(11), Z =>
                           mult_143_n6203);
   mult_143_U4644 : XOR2_X1 port map( A => n3718, B => n3681, Z => n1665);
   mult_143_U4640 : XOR2_X1 port map( A => mult_143_n6192, B => A_SIG(8), Z => 
                           n1663);
   mult_143_U4639 : XOR2_X1 port map( A => mult_143_n6189, B => A_SIG(11), Z =>
                           n1662);
   mult_143_U4638 : XOR2_X1 port map( A => n3717, B => n3716, Z => 
                           mult_143_n6186);
   mult_143_U4637 : XOR2_X1 port map( A => n649, B => mult_143_n6184, Z => 
                           mult_143_n6168);
   mult_143_U4635 : XOR2_X1 port map( A => mult_143_n6170, B => A_SIG(11), Z =>
                           n1661);
   mult_143_U4634 : XOR2_X1 port map( A => mult_143_n6165, B => A_SIG(8), Z => 
                           n1660);
   mult_143_U4633 : XOR2_X1 port map( A => n3714, B => n3680, Z => 
                           mult_143_n6162);
   mult_143_U4632 : XOR2_X1 port map( A => mult_143_n6158, B => A_SIG(11), Z =>
                           mult_143_n6148);
   mult_143_U4631 : XOR2_X1 port map( A => A_SIG(11), B => mult_143_n6157, Z =>
                           mult_143_n6147);
   mult_143_U4630 : XOR2_X1 port map( A => mult_143_n6154, B => A_SIG(11), Z =>
                           n1659);
   mult_143_U4626 : XOR2_X1 port map( A => mult_143_n6143, B => A_SIG(8), Z => 
                           mult_143_n6137);
   mult_143_U4625 : XOR2_X1 port map( A => A_SIG(8), B => mult_143_n6142, Z => 
                           mult_143_n6136);
   mult_143_U4624 : XOR2_X1 port map( A => mult_143_n6139, B => A_SIG(8), Z => 
                           mult_143_n5412);
   mult_143_U4621 : XOR2_X1 port map( A => n642, B => mult_143_n6132, Z => 
                           mult_143_n5128);
   mult_143_U4580 : XOR2_X1 port map( A => n3774, B => n3581, Z => n1657);
   mult_143_U4575 : XOR2_X1 port map( A => mult_143_n5960, B => n3793, Z => 
                           n1039);
   mult_143_U4517 : XOR2_X1 port map( A => n4634, B => n2617, Z => 
                           mult_143_n5794);
   mult_143_U4516 : XOR2_X1 port map( A => mult_143_n1893, B => n2630, Z => 
                           mult_143_n5793);
   mult_143_U4515 : XOR2_X1 port map( A => n3796, B => n3061, Z => 
                           mult_143_n5783);
   mult_143_U4514 : XOR2_X1 port map( A => mult_143_n5780, B => mult_143_n5781,
                           Z => mult_143_n5779);
   mult_143_U4511 : XOR2_X1 port map( A => mult_143_n5768, B => mult_143_n5758,
                           Z => n1650);
   mult_143_U4501 : XOR2_X1 port map( A => n2714, B => mult_143_n5531, Z => 
                           mult_143_n5755);
   mult_143_U4500 : XOR2_X1 port map( A => n2692, B => mult_143_n5755, Z => 
                           n1649);
   mult_143_U4499 : XOR2_X1 port map( A => mult_143_n5754, B => n3709, Z => 
                           mult_143_n5435);
   mult_143_U4491 : XOR2_X1 port map( A => n2665, B => n3058, Z => 
                           mult_143_n5746);
   mult_143_U4489 : XOR2_X1 port map( A => mult_143_n5742, B => mult_143_n5743,
                           Z => mult_143_n5740);
   mult_143_U4478 : XOR2_X1 port map( A => n4586, B => n3803, Z => 
                           mult_143_n5686);
   mult_143_U4477 : XOR2_X1 port map( A => n3067, B => n2747, Z => 
                           mult_143_n5693);
   mult_143_U4476 : XOR2_X1 port map( A => mult_143_n2759, B => mult_143_n6367,
                           Z => mult_143_n5692);
   mult_143_U4475 : XOR2_X1 port map( A => n4689, B => mult_143_n5686, Z => 
                           mult_143_n5684);
   mult_143_U4472 : XOR2_X1 port map( A => mult_143_n6590, B => n1628, Z => 
                           mult_143_n5673);
   mult_143_U4471 : XOR2_X1 port map( A => n4585, B => n2750, Z => 
                           mult_143_n5672);
   mult_143_U4468 : XOR2_X1 port map( A => mult_143_n6583, B => n4946, Z => 
                           mult_143_n5657);
   mult_143_U4467 : XOR2_X1 port map( A => mult_143_n5656, B => mult_143_n5657,
                           Z => n1643);
   mult_143_U4464 : XOR2_X1 port map( A => mult_143_n5632, B => mult_143_n5228,
                           Z => mult_143_n5597);
   mult_143_U4463 : XOR2_X1 port map( A => mult_143_n5628, B => mult_143_n5619,
                           Z => mult_143_n5615);
   mult_143_U4462 : XOR2_X1 port map( A => n3632, B => n3628, Z => 
                           mult_143_n5622);
   mult_143_U4461 : XOR2_X1 port map( A => mult_143_n5612, B => n2759, Z => 
                           mult_143_n5620);
   mult_143_U4460 : XOR2_X1 port map( A => mult_143_n6541, B => n2615, Z => 
                           mult_143_n5618);
   mult_143_U4459 : XOR2_X1 port map( A => mult_143_n5418, B => mult_143_n5618,
                           Z => mult_143_n5425);
   mult_143_U4457 : XOR2_X1 port map( A => mult_143_n5425, B => n4764, Z => 
                           mult_143_n5614);
   mult_143_U4454 : XOR2_X1 port map( A => mult_143_n5419, B => mult_143_n5420,
                           Z => mult_143_n5609);
   mult_143_U4449 : XOR2_X1 port map( A => mult_143_n5598, B => mult_143_n5597,
                           Z => mult_143_n5595);
   mult_143_U4446 : XOR2_X1 port map( A => n2859, B => mult_143_n5585, Z => 
                           mult_143_n5215);
   mult_143_U4445 : XOR2_X1 port map( A => mult_143_n5582, B => mult_143_n5583,
                           Z => mult_143_n5581);
   mult_143_U4443 : XOR2_X1 port map( A => n3633, B => n3626, Z => 
                           mult_143_n5567);
   mult_143_U4439 : XOR2_X1 port map( A => mult_143_n6402, B => mult_143_n5564,
                           Z => mult_143_n5563);
   mult_143_U4438 : XOR2_X1 port map( A => mult_143_n5562, B => mult_143_n5563,
                           Z => mult_143_n5396);
   mult_143_U4433 : XOR2_X1 port map( A => mult_143_n6417, B => n4575, Z => 
                           mult_143_n5550);
   mult_143_U4431 : XOR2_X1 port map( A => mult_143_n5542, B => mult_143_n5543,
                           Z => mult_143_n5541);
   mult_143_U4430 : XOR2_X1 port map( A => n2726, B => n3795, Z => 
                           mult_143_n5539);
   mult_143_U4429 : XOR2_X1 port map( A => n3050, B => mult_143_n5539, Z => 
                           n1640);
   mult_143_U4428 : XOR2_X1 port map( A => mult_143_n6322, B => mult_143_n5527,
                           Z => mult_143_n5526);
   mult_143_U4427 : XOR2_X1 port map( A => mult_143_n5525, B => mult_143_n5526,
                           Z => n1639);
   mult_143_U4419 : XOR2_X1 port map( A => mult_143_n5524, B => mult_143_n5523,
                           Z => mult_143_n5522);
   mult_143_U4411 : XOR2_X1 port map( A => mult_143_n5517, B => n3700, Z => 
                           mult_143_n5221);
   mult_143_U4409 : XOR2_X1 port map( A => mult_143_n5495, B => n3591, Z => 
                           mult_143_n5485);
   mult_143_U4408 : XOR2_X1 port map( A => A_SIG(17), B => mult_143_n5489, Z =>
                           n1637);
   mult_143_U4407 : XOR2_X1 port map( A => A_SIG(20), B => mult_143_n5486, Z =>
                           n1636);
   mult_143_U4401 : XOR2_X1 port map( A => mult_143_n5461, B => n2715, Z => 
                           n1635);
   mult_143_U4400 : XOR2_X1 port map( A => n3707, B => n3818, Z => 
                           mult_143_n5450);
   mult_143_U4392 : XOR2_X1 port map( A => n748, B => mult_143_n5403, Z => 
                           mult_143_n4850);
   mult_143_U4391 : XOR2_X1 port map( A => n748, B => mult_143_n5402, Z => 
                           mult_143_n4831);
   mult_143_U4388 : XOR2_X1 port map( A => n962, B => mult_143_n5381, Z => 
                           mult_143_n5379);
   mult_143_U4384 : XOR2_X1 port map( A => mult_143_n6479, B => mult_143_n6478,
                           Z => mult_143_n5362);
   mult_143_U4383 : XOR2_X1 port map( A => n2632, B => n4588, Z => 
                           mult_143_n5361);
   mult_143_U4371 : XOR2_X1 port map( A => mult_143_n5329, B => n2612, Z => 
                           mult_143_n5288);
   mult_143_U4367 : XOR2_X1 port map( A => mult_143_n5272, B => n2723, Z => 
                           mult_143_n5270);
   mult_143_U4360 : XOR2_X1 port map( A => n4750, B => n3547, Z => n1632);
   mult_143_U4351 : XOR2_X1 port map( A => mult_143_n5138, B => mult_143_n5137,
                           Z => mult_143_n5132);
   mult_143_U4349 : XOR2_X1 port map( A => n536, B => mult_143_n5134, Z => 
                           mult_143_n5133);
   mult_143_U4348 : XOR2_X1 port map( A => n536, B => mult_143_n5129, Z => 
                           mult_143_n5117);
   mult_143_U4347 : XOR2_X1 port map( A => mult_143_n5127, B => mult_143_n5128,
                           Z => mult_143_n5118);
   mult_143_U4339 : MUX2_X1 port map( A => n3795, B => n4634, S => n2780, Z => 
                           mult_143_n610);
   mult_143_U4332 : XOR2_X1 port map( A => n4634, B => mult_143_n1897, Z => 
                           mult_143_n5095);
   mult_143_U4327 : XOR2_X1 port map( A => mult_143_n1816, B => mult_143_n5074,
                           Z => n1630);
   mult_143_U4316 : XOR2_X1 port map( A => n1560, B => n4768, Z => 
                           mult_143_n5020);
   mult_143_U4312 : XOR2_X1 port map( A => n2840, B => mult_143_n5007, Z => 
                           n1628);
   mult_143_U4309 : XOR2_X1 port map( A => n3775, B => n3551, Z => 
                           mult_143_n4994);
   mult_143_U4301 : XOR2_X1 port map( A => n4760, B => n3541, Z => 
                           mult_143_n4965);
   mult_143_U4300 : XOR2_X1 port map( A => n3504, B => n4590, Z => 
                           mult_143_n4966);
   mult_143_U4294 : XOR2_X1 port map( A => n4630, B => n4590, Z => 
                           mult_143_n4949);
   mult_143_U4291 : XOR2_X1 port map( A => n3797, B => n3565, Z => n1627);
   mult_143_U4290 : XOR2_X1 port map( A => n3775, B => n3563, Z => n1626);
   mult_143_U4288 : XOR2_X1 port map( A => n4760, B => mult_143_n4925, Z => 
                           n1625);
   mult_143_U4287 : XOR2_X1 port map( A => n4750, B => mult_143_n4922, Z => 
                           n1624);
   mult_143_U4283 : XOR2_X1 port map( A => n1572, B => n4630, Z => 
                           mult_143_n4897);
   mult_143_U4282 : XOR2_X1 port map( A => n3796, B => n3570, Z => n1623);
   mult_143_U4281 : XOR2_X1 port map( A => n748, B => mult_143_n4889, Z => 
                           n1622);
   mult_143_U4279 : XOR2_X1 port map( A => n3691, B => n1621, Z => 
                           mult_143_n4883);
   mult_143_U4278 : XOR2_X1 port map( A => n4760, B => n3545, Z => n1620);
   mult_143_U4277 : XOR2_X1 port map( A => n1613, B => n1620, Z => 
                           mult_143_n4870);
   mult_143_U4273 : XOR2_X1 port map( A => n1590, B => n1614, Z => 
                           mult_143_n4853);
   mult_143_U4271 : XOR2_X1 port map( A => mult_143_n4846, B => A_SIG(8), Z => 
                           n1618);
   mult_143_U4269 : XOR2_X1 port map( A => n3568, B => n3794, Z => n1617);
   mult_143_U4268 : XOR2_X1 port map( A => A_SIG(17), B => mult_143_n4822, Z =>
                           n1616);
   mult_143_U4267 : XOR2_X1 port map( A => n3689, B => n3651, Z => 
                           mult_143_n4815);
   mult_143_U4266 : XOR2_X1 port map( A => n2614, B => mult_143_n4807, Z => 
                           SIG_in(3));
   mult_143_U4265 : XOR2_X1 port map( A => n963, B => n2602, Z => SIG_in(6));
   mult_143_U4264 : XOR2_X1 port map( A => mult_143_n4798, B => mult_143_n4799,
                           Z => SIG_in(9));
   mult_143_U4263 : XOR2_X1 port map( A => mult_143_n4797, B => n4697, Z => 
                           SIG_in(10));
   mult_143_U4262 : NAND3_X1 port map( A1 => n4697, A2 => mult_143_n4401, A3 =>
                           n4901, ZN => mult_143_n4791);
   mult_143_U4261 : XOR2_X1 port map( A => mult_143_n4793, B => mult_143_n4794,
                           Z => SIG_in(12));
   mult_143_U4260 : XOR2_X1 port map( A => n2637, B => mult_143_n4790, Z => 
                           SIG_in(13));
   mult_143_U4259 : XOR2_X1 port map( A => n720, B => mult_143_n4786, Z => 
                           SIG_in(14));
   mult_143_U4258 : XOR2_X1 port map( A => n4756, B => mult_143_n4783, Z => 
                           SIG_in(16));
   mult_143_U4257 : XOR2_X1 port map( A => mult_143_n4778, B => mult_143_n4779,
                           Z => SIG_in(18));
   mult_143_U4256 : XOR2_X1 port map( A => n3642, B => n3577, Z => SIG_in(19));
   mult_143_U4255 : XOR2_X1 port map( A => n3828, B => n3743, Z => SIG_in(20));
   mult_143_U4254 : XOR2_X1 port map( A => n3614, B => n1541, Z => SIG_in(22));
   mult_143_U4027 : MUX2_X1 port map( A => mult_143_n4555, B => n630, S => 
                           B_SIG(2), Z => mult_143_n6230);
   mult_143_U3783 : OAI21_X1 port map( B1 => n3643, B2 => n1589, A => 
                           mult_143_n1942, ZN => n1531);
   mult_143_U3714 : OAI21_X1 port map( B1 => n3645, B2 => n1589, A => 
                           mult_143_n2001, ZN => mult_143_n6067);
   mult_143_U3597 : AOI21_X1 port map( B1 => n4890, B2 => n4664, A => 
                           mult_143_n5997, ZN => n1530);
   mult_143_U3586 : OAI21_X1 port map( B1 => n3644, B2 => n1589, A => 
                           mult_143_n2200, ZN => mult_143_n5986);
   mult_143_U3511 : OAI21_X1 port map( B1 => n3597, B2 => n1589, A => n3517, ZN
                           => n1529);
   mult_143_U3447 : OAI21_X1 port map( B1 => n3659, B2 => n1589, A => 
                           mult_143_n2401, ZN => mult_143_n5855);
   mult_143_U3302 : AOI21_X1 port map( B1 => mult_143_n6570, B2 => n3067, A => 
                           n3803, ZN => mult_143_n5735);
   mult_143_U3301 : NOR2_X1 port map( A1 => n3067, A2 => mult_143_n6570, ZN => 
                           mult_143_n5736);
   mult_143_U3255 : AOI22_X1 port map( A1 => mult_143_n6605, A2 => n4657, B1 =>
                           n3803, B2 => n955, ZN => mult_143_n5691);
   mult_143_U3254 : XNOR2_X1 port map( A => n2707, B => mult_143_n5691, ZN => 
                           mult_143_n5652);
   mult_143_U3007 : NAND2_X1 port map( A1 => mult_143_n4991, A2 => n2864, ZN =>
                           mult_143_n2759);
   mult_143_U2843 : AOI21_X1 port map( B1 => mult_143_n5232, B2 => n3503, A => 
                           mult_143_n426, ZN => mult_143_n5236);
   mult_143_U2805 : NOR2_X1 port map( A1 => mult_143_n5189, A2 => 
                           mult_143_n5190, ZN => n949);
   mult_143_U2804 : AOI21_X1 port map( B1 => mult_143_n5187, B2 => n4763, A => 
                           n949, ZN => n1055);
   mult_143_U2578 : AOI222_X1 port map( A1 => mult_143_n4956, A2 => n657, B1 =>
                           mult_143_n4956, B2 => mult_143_n6367, C1 => n657, C2
                           => mult_143_n6367, ZN => mult_143_n813);
   mult_143_U2552 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => 
                           mult_143_n4891, A => mult_143_n4933, ZN => 
                           mult_143_n4932);
   mult_143_U2551 : AOI21_X1 port map( B1 => B_SIG(7), B2 => mult_143_n96, A =>
                           mult_143_n4932, ZN => mult_143_n4931);
   mult_143_n4468 <= '0';
   mult_143_n4467 <= '1';
   mult_143_n4327 <= '0';
   mult_143_n4325 <= '0';
   mult_143_n4319 <= '0';
   mult_143_n4317 <= '0';
   mult_143_n4309 <= '0';
   mult_143_n4307 <= '0';
   mult_143_n4301 <= '0';
   mult_143_n4275 <= '0';
   mult_143_n4273 <= '0';
   mult_143_n4217 <= '0';
   mult_143_n4215 <= '0';
   mult_143_n4208 <= '0';
   mult_143_n4206 <= '0';
   mult_143_n4201 <= '0';
   mult_143_n4199 <= '0';
   mult_143_n4156 <= '0';
   mult_143_n4154 <= '0';
   mult_143_MY_CLK_r_REG423_S1 : DFF_X1 port map( D => mult_143_n655, CK => clk
                           , Q => n_1168, QN => mult_143_n6346);
   mult_143_MY_CLK_r_REG422_S1 : DFF_X1 port map( D => mult_143_n654, CK => clk
                           , Q => n_1169, QN => mult_143_n6582);
   mult_143_U2618 : XNOR2_X1 port map( A => mult_143_n4994, B => mult_143_n4995
                           , ZN => mult_143_n6597);
   mult_143_U3001 : AOI21_X1 port map( B1 => n2918, B2 => mult_143_n5430, A => 
                           mult_143_n5431, ZN => mult_143_n276);
   mult_143_U2894 : XNOR2_X1 port map( A => n1740, B => n1739, ZN => 
                           mult_143_n5318);
   mult_143_U2914 : XNOR2_X1 port map( A => mult_143_n5276, B => mult_143_n5275
                           , ZN => mult_143_n5338);
   mult_143_U2676 : OAI21_X1 port map( B1 => n3655, B2 => n3643, A => 
                           mult_143_n5047, ZN => mult_143_n5046);
   mult_143_U2890 : XNOR2_X1 port map( A => n3622, B => n3612, ZN => 
                           mult_143_n5315);
   mult_143_U2569 : XNOR2_X1 port map( A => mult_143_n4948, B => mult_143_n4949
                           , ZN => n964);
   mult_143_U2922 : XNOR2_X1 port map( A => n2865, B => n3091, ZN => 
                           mult_143_n5342);
   mult_143_U3653 : NOR2_X1 port map( A1 => mult_143_n6028, A2 => n865, ZN => 
                           mult_143_n6027);
   mult_143_U2485 : XNOR2_X1 port map( A => mult_143_n4862, B => n4754, ZN => 
                           n1614);
   mult_143_U2808 : NOR2_X1 port map( A1 => n1632, A2 => n1588, ZN => 
                           mult_143_n4344);
   mult_143_U2806 : OAI21_X1 port map( B1 => n3099, B2 => n4670, A => 
                           mult_143_n5191, ZN => n991);
   mult_143_U2590 : XNOR2_X1 port map( A => mult_143_n4965, B => mult_143_n4966
                           , ZN => mult_143_n812);
   mult_143_U3651 : AOI22_X1 port map( A1 => mult_143_n6027, A2 => n868, B1 => 
                           mult_143_n6028, B2 => n865, ZN => mult_143_n6026);
   mult_143_U2609 : AOI21_X1 port map( B1 => n4736, B2 => n3806, A => 
                           mult_143_n4987, ZN => n1528);
   mult_143_U2490 : XNOR2_X1 port map( A => mult_143_n4870, B => mult_143_n4869
                           , ZN => n968);
   mult_143_U2500 : XNOR2_X1 port map( A => mult_143_n4490, B => mult_143_n4879
                           , ZN => n1613);
   mult_143_U2918 : XNOR2_X1 port map( A => n3634, B => n4615, ZN => 
                           mult_143_n5340);
   mult_143_U2828 : XNOR2_X1 port map( A => n1633, B => n1561, ZN => 
                           mult_143_n5142);
   mult_143_U3676 : XNOR2_X1 port map( A => n4760, B => mult_143_n6043, ZN => 
                           mult_143_n1610);
   mult_143_U2703 : AOI21_X1 port map( B1 => n2908, B2 => n3806, A => 
                           mult_143_n5070, ZN => mult_143_n5069);
   mult_143_U2967 : AOI21_X1 port map( B1 => n3510, B2 => n3742, A => n1698, ZN
                           => mult_143_n6620);
   U19 : NAND2_X1 port map( A1 => n378, A2 => n544, ZN => n542);
   U20 : NAND2_X1 port map( A1 => mult_143_n5299, A2 => n1048, ZN => n378);
   U23 : NAND2_X1 port map( A1 => mult_143_n5012, A2 => n381, ZN => n380);
   U24 : NAND2_X1 port map( A1 => n772, A2 => B_SIG(19), ZN => n381);
   U48 : AND2_X1 port map( A1 => mult_143_n5263, A2 => mult_143_n5264, ZN => 
                           n386);
   U52 : NAND2_X1 port map( A1 => n1488, A2 => n1047, ZN => n388);
   U55 : NAND2_X1 port map( A1 => mult_143_n5350, A2 => n392, ZN => n391);
   U56 : NAND2_X1 port map( A1 => mult_143_n6532, A2 => n2713, ZN => n392);
   U65 : NOR2_X1 port map( A1 => B_SIG(11), A2 => n2841, ZN => n398);
   U67 : NAND2_X1 port map( A1 => B_SIG(11), A2 => n2841, ZN => n400);
   U71 : NAND2_X1 port map( A1 => mult_143_n6109, A2 => n404, ZN => n403);
   U72 : NAND2_X1 port map( A1 => n3820, A2 => n3804, ZN => n404);
   U77 : NAND2_X1 port map( A1 => n3806, A2 => n3804, ZN => n408);
   U89 : AOI21_X1 port map( B1 => mult_143_n2755, B2 => mult_143_n5434, A => 
                           mult_143_n5435, ZN => n512);
   U91 : OR2_X1 port map( A1 => mult_143_n5582, A2 => mult_143_n5583, ZN => 
                           n416);
   U92 : AND2_X1 port map( A1 => mult_143_n5582, A2 => mult_143_n5583, ZN => 
                           n417);
   U95 : NAND2_X1 port map( A1 => n420, A2 => n419, ZN => n418);
   U97 : INV_X1 port map( A => mult_143_n5594, ZN => n420);
   U98 : NAND2_X1 port map( A1 => n422, A2 => mult_143_n5631, ZN => n421);
   U99 : NAND2_X1 port map( A1 => mult_143_n5594, A2 => mult_143_n6607, ZN => 
                           n422);
   U102 : NAND2_X1 port map( A1 => n426, A2 => n425, ZN => n424);
   U114 : OAI21_X1 port map( B1 => n3613, B2 => n3645, A => n434, ZN => n433);
   U116 : INV_X1 port map( A => mult_143_n5065, ZN => n435);
   U123 : NAND2_X1 port map( A1 => n2825, A2 => mult_143_n6002, ZN => n440);
   U133 : AND2_X1 port map( A1 => n3817, A2 => n4695, ZN => n446);
   U146 : NAND2_X1 port map( A1 => mult_143_n867, A2 => n1040, ZN => n453);
   U149 : NAND2_X1 port map( A1 => mult_143_n5057, A2 => n457, ZN => n456);
   U150 : NAND2_X1 port map( A1 => mult_143_n72, A2 => B_SIG(20), ZN => n457);
   U160 : OR2_X1 port map( A1 => mult_143_n5730, A2 => mult_143_n5731, ZN => 
                           n463);
   U161 : AND2_X1 port map( A1 => mult_143_n5730, A2 => mult_143_n5731, ZN => 
                           n464);
   U164 : NAND3_X1 port map( A1 => mult_143_n6287, A2 => n809, A3 => n808, ZN 
                           => n812);
   U166 : MUX2_X1 port map( A => n4580, B => n3588, S => n1567, Z => 
                           mult_143_n4995);
   U177 : XNOR2_X1 port map( A => n3748, B => n4610, ZN => n473);
   U185 : INV_X1 port map( A => mult_143_n6104, ZN => n479);
   U192 : NOR2_X1 port map( A1 => n485, A2 => n484, ZN => mult_143_n5489);
   U193 : INV_X1 port map( A => mult_143_n5491, ZN => n484);
   U200 : AND3_X1 port map( A1 => mult_143_n6287, A2 => n809, A3 => n808, ZN =>
                           n825);
   U201 : NAND2_X1 port map( A1 => n891, A2 => B_SIG(8), ZN => n490);
   U216 : NAND2_X1 port map( A1 => mult_143_n5054, A2 => n501, ZN => n500);
   U217 : NAND2_X1 port map( A1 => n3806, A2 => n4695, ZN => n501);
   U228 : XNOR2_X1 port map( A => mult_143_n5092, B => n1839, ZN => 
                           mult_143_n5086);
   U237 : OR2_X1 port map( A1 => mult_143_n5465, A2 => mult_143_n5466, ZN => 
                           n513);
   U240 : NAND2_X1 port map( A1 => n518, A2 => n3602, ZN => n516);
   U242 : NAND2_X1 port map( A1 => n1520, A2 => n3502, ZN => n518);
   U243 : OR2_X1 port map( A1 => n4851, A2 => n3502, ZN => n519);
   U260 : NOR2_X1 port map( A1 => n637, A2 => n587, ZN => mult_143_n6097);
   U263 : MUX2_X1 port map( A => mult_143_n6367, B => n4730, S => n657, Z => 
                           mult_143_n4957);
   U272 : NAND2_X1 port map( A1 => n878, A2 => B_SIG(9), ZN => n539);
   U276 : NAND2_X1 port map( A1 => n542, A2 => n821, ZN => mult_143_n5284);
   U281 : XNOR2_X1 port map( A => mult_143_n5672, B => n3831, ZN => 
                           mult_143_n5667);
   U284 : OR2_X1 port map( A1 => n1562, A2 => n3706, ZN => n547);
   U285 : AND2_X1 port map( A1 => n1562, A2 => n3706, ZN => n548);
   U286 : OAI21_X1 port map( B1 => mult_143_n5646, B2 => n552, A => n549, ZN =>
                           mult_143_n5671);
   U287 : NAND2_X1 port map( A1 => n4642, A2 => n3138, ZN => n549);
   U290 : AND2_X1 port map( A1 => mult_143_n5648, A2 => mult_143_n5647, ZN => 
                           n552);
   U297 : OAI21_X1 port map( B1 => mult_143_n6113, B2 => B_SIG(21), A => 
                           B_SIG(22), ZN => mult_143_n6114);
   U312 : AND2_X1 port map( A1 => mult_143_n5722, A2 => mult_143_n5723, ZN => 
                           n563);
   U313 : NAND3_X1 port map( A1 => n1070, A2 => n809, A3 => n808, ZN => 
                           mult_143_n6079);
   U316 : NAND2_X1 port map( A1 => mult_143_n4849, A2 => n565, ZN => n564);
   U317 : NAND2_X1 port map( A1 => mult_143_n36, A2 => B_SIG(14), ZN => n565);
   U318 : INV_X1 port map( A => mult_143_n4848, ZN => n566);
   U319 : INV_X1 port map( A => mult_143_n6625, ZN => n567);
   U321 : AND2_X1 port map( A1 => n4675, A2 => n3806, ZN => n569);
   U325 : AND2_X1 port map( A1 => n1027, A2 => B_SIG(16), ZN => n572);
   U326 : INV_X1 port map( A => mult_143_n6124, ZN => n573);
   U327 : NAND2_X1 port map( A1 => n573, A2 => n1077, ZN => n826);
   U328 : XNOR2_X1 port map( A => mult_143_n5999, B => n852, ZN => n1557);
   U339 : NAND2_X1 port map( A1 => n584, A2 => n581, ZN => mult_143_n5268);
   U345 : INV_X1 port map( A => mult_143_n6041, ZN => n585);
   U347 : NAND2_X1 port map( A1 => n573, A2 => n1032, ZN => n587);
   U362 : NAND2_X1 port map( A1 => n1032, A2 => mult_143_n6118, ZN => n599);
   U373 : OAI22_X1 port map( A1 => mult_143_n6095, A2 => B_SIG(19), B1 => 
                           mult_143_n6040, B2 => mult_143_n6096, ZN => n607);
   U376 : NAND2_X1 port map( A1 => n611, A2 => n4571, ZN => n813);
   U378 : NAND2_X1 port map( A1 => mult_143_n5232, A2 => mult_143_n427, ZN => 
                           n611);
   U385 : NAND2_X1 port map( A1 => mult_143_n6397, A2 => mult_143_n6398, ZN => 
                           n616);
   U388 : AOI21_X1 port map( B1 => n624, B2 => n2786, A => mult_143_n6578, ZN 
                           => mult_143_n4761);
   U389 : AOI21_X1 port map( B1 => mult_143_n4759, B2 => n2784, A => 
                           mult_143_n6560, ZN => mult_143_n4757);
   U409 : INV_X1 port map( A => mult_143_n5732, ZN => n716);
   U413 : INV_X1 port map( A => mult_143_n5671, ZN => n1836);
   U420 : INV_X1 port map( A => mult_143_n3448, ZN => n743);
   U421 : INV_X1 port map( A => n4882, ZN => n744);
   U432 : NAND2_X1 port map( A1 => mult_143_n6079, A2 => mult_143_n6260, ZN => 
                           mult_143_n6126);
   U433 : INV_X1 port map( A => mult_143_n6036, ZN => n637);
   U434 : AOI22_X1 port map( A1 => n637, A2 => n860, B1 => B_SIG(16), B2 => 
                           n2906, ZN => mult_143_n6035);
   U435 : OAI21_X1 port map( B1 => n3647, B2 => n3644, A => mult_143_n4946, ZN 
                           => mult_143_n4945);
   U436 : OAI21_X1 port map( B1 => n3647, B2 => n3596, A => mult_143_n5041, ZN 
                           => mult_143_n5040);
   U438 : OAI21_X1 port map( B1 => n3647, B2 => n3673, A => mult_143_n4902, ZN 
                           => mult_143_n4901);
   U439 : OAI21_X1 port map( B1 => n3647, B2 => n3643, A => mult_143_n6093, ZN 
                           => mult_143_n6092);
   U440 : OAI21_X1 port map( B1 => n3647, B2 => n3597, A => mult_143_n5907, ZN 
                           => mult_143_n5906);
   U441 : OAI21_X1 port map( B1 => n3647, B2 => n3659, A => mult_143_n5846, ZN 
                           => mult_143_n5845);
   U442 : OAI21_X1 port map( B1 => n3647, B2 => n3594, A => n1498, ZN => 
                           mult_143_n6005);
   U443 : OAI21_X1 port map( B1 => B_SIG(3), B2 => B_SIG(4), A => n2823, ZN => 
                           mult_143_n6289);
   U444 : AOI221_X1 port map( B1 => B_SIG(3), B2 => B_SIG(4), C1 => 
                           mult_143_n6290, C2 => B_SIG(4), A => B_SIG(5), ZN =>
                           mult_143_n6286);
   U446 : OAI21_X1 port map( B1 => n3687, B2 => n3673, A => mult_143_n5949, ZN 
                           => mult_143_n5948);
   U447 : OAI21_X1 port map( B1 => n1557, B2 => mult_143_n5859, A => 
                           mult_143_n5901, ZN => mult_143_n5900);
   U448 : OAI21_X1 port map( B1 => n1557, B2 => mult_143_n4828, A => 
                           mult_143_n5982, ZN => mult_143_n5981);
   U450 : OAI21_X1 port map( B1 => n3649, B2 => n3594, A => mult_143_n5998, ZN 
                           => mult_143_n5997);
   U451 : XNOR2_X1 port map( A => n3776, B => n3744, ZN => SIG_in(26));
   U452 : NAND2_X1 port map( A1 => mult_143_n6289, A2 => mult_143_n6288, ZN => 
                           mult_143_n6272);
   U453 : NAND2_X1 port map( A1 => n1069, A2 => mult_143_n6127, ZN => 
                           mult_143_n6022);
   U455 : OAI21_X1 port map( B1 => n3640, B2 => mult_143_n5306, A => 
                           mult_143_n5307, ZN => mult_143_n5303);
   U456 : AND2_X1 port map( A1 => mult_143_n5268, A2 => mult_143_n5269, ZN => 
                           mult_143_n5271);
   U457 : OAI22_X1 port map( A1 => mult_143_n5268, A2 => mult_143_n5269, B1 => 
                           mult_143_n5271, B2 => mult_143_n5270, ZN => 
                           mult_143_n5256);
   U458 : OAI221_X1 port map( B1 => mult_143_n430, B2 => mult_143_n6620, C1 => 
                           mult_143_n6619, C2 => n2890, A => mult_143_n5236, ZN
                           => mult_143_n5235);
   U459 : OAI21_X1 port map( B1 => n3654, B2 => n3596, A => mult_143_n6045, ZN 
                           => n1527);
   U460 : OAI21_X1 port map( B1 => n3654, B2 => n3673, A => mult_143_n5958, ZN 
                           => n1526);
   U461 : OAI21_X1 port map( B1 => n3654, B2 => n3597, A => mult_143_n5913, ZN 
                           => mult_143_n5912);
   U462 : OAI21_X1 port map( B1 => n3654, B2 => n3659, A => mult_143_n5852, ZN 
                           => n1525);
   U463 : XNOR2_X1 port map( A => mult_143_n4972, B => mult_143_n4973, ZN => 
                           n994);
   U464 : XNOR2_X1 port map( A => n817, B => mult_143_n4760, ZN => SIG_in(24));
   U467 : NAND2_X1 port map( A1 => mult_143_n4788, A2 => mult_143_n4791, ZN => 
                           mult_143_n4794);
   U468 : OAI21_X1 port map( B1 => n3676, B2 => n3594, A => mult_143_n5200, ZN 
                           => mult_143_n5199);
   U469 : OAI21_X1 port map( B1 => n3676, B2 => n3643, A => mult_143_n6101, ZN 
                           => mult_143_n6100);
   U470 : OAI21_X1 port map( B1 => n3676, B2 => n3645, A => mult_143_n6065, ZN 
                           => mult_143_n6064);
   U471 : OAI21_X1 port map( B1 => mult_143_n4407, B2 => mult_143_n4848, A => 
                           mult_143_n5955, ZN => n1524);
   U473 : OAI21_X1 port map( B1 => n3676, B2 => n3644, A => mult_143_n5985, ZN 
                           => mult_143_n5984);
   U474 : OAI21_X1 port map( B1 => n3676, B2 => n3659, A => mult_143_n5849, ZN 
                           => n1523);
   U480 : OAI21_X1 port map( B1 => n3613, B2 => n3597, A => mult_143_n5904, ZN 
                           => mult_143_n5903);
   U481 : OAI21_X1 port map( B1 => n1024, B2 => mult_143_n4824, A => 
                           mult_143_n6039, ZN => mult_143_n6038);
   U482 : OAI21_X1 port map( B1 => n3613, B2 => n3673, A => mult_143_n5952, ZN 
                           => mult_143_n5951);
   U485 : OR2_X1 port map( A1 => mult_143_n6286, A2 => n895, ZN => n809);
   U487 : AOI21_X1 port map( B1 => n826, B2 => mult_143_n6002, A => 
                           mult_143_n6003, ZN => mult_143_n6000);
   U489 : AOI22_X1 port map( A1 => B_SIG(1), A2 => mult_143_n74, B1 => 
                           mult_143_n76, B2 => B_SIG(0), ZN => mult_143_n6295);
   U490 : AOI22_X1 port map( A1 => mult_143_n74, A2 => B_SIG(2), B1 => 
                           mult_143_n84, B2 => B_SIG(0), ZN => mult_143_n6299);
   U491 : AOI22_X1 port map( A1 => B_SIG(2), A2 => n2598, B1 => B_SIG(0), B2 =>
                           mult_143_n96, ZN => mult_143_n5405);
   U492 : AOI22_X1 port map( A1 => B_SIG(2), A2 => n765, B1 => B_SIG(0), B2 => 
                           mult_143_n48, ZN => mult_143_n6160);
   U493 : AOI221_X1 port map( B1 => B_SIG(1), B2 => n774, C1 => B_SIG(0), C2 =>
                           mult_143_n72, A => mult_143_n6234, ZN => 
                           mult_143_n6233);
   U494 : AOI221_X1 port map( B1 => n804, B2 => B_SIG(1), C1 => B_SIG(0), C2 =>
                           mult_143_n6621, A => mult_143_n6183, ZN => 
                           mult_143_n6182);
   U495 : AOI22_X1 port map( A1 => B_SIG(2), A2 => n755, B1 => B_SIG(0), B2 => 
                           mult_143_n36, ZN => mult_143_n6145);
   U496 : NAND2_X1 port map( A1 => B_SIG(0), A2 => n651, ZN => n1612);
   U497 : AOI21_X1 port map( B1 => B_SIG(0), B2 => n646, A => n1765, ZN => 
                           mult_143_n6146);
   U498 : AOI221_X1 port map( B1 => n1031, B2 => B_SIG(1), C1 => B_SIG(0), C2 
                           => mult_143_n3228, A => mult_143_n6134, ZN => 
                           mult_143_n6133);
   U499 : NAND2_X1 port map( A1 => B_SIG(0), A2 => n748, ZN => mult_143_n2743);
   U500 : NAND2_X1 port map( A1 => B_SIG(0), A2 => n650, ZN => n1611);
   U501 : NAND2_X1 port map( A1 => B_SIG(0), A2 => n646, ZN => mult_143_n5413);
   U502 : NAND2_X1 port map( A1 => B_SIG(0), A2 => n648, ZN => n1610);
   U503 : NOR2_X1 port map( A1 => mult_143_n4945, A2 => n811, ZN => 
                           mult_143_n4944);
   U506 : OAI21_X1 port map( B1 => n874, B2 => n882, A => n878, ZN => 
                           mult_143_n6259);
   U508 : AOI21_X1 port map( B1 => n874, B2 => n882, A => n878, ZN => 
                           mult_143_n6258);
   U514 : OR2_X1 port map( A1 => mult_143_n427, A2 => mult_143_n5232, ZN => 
                           n814);
   U517 : OAI21_X1 port map( B1 => B_SIG(22), B2 => mult_143_n6113, A => 
                           mult_143_n6114, ZN => mult_143_n6112);
   U519 : INV_X1 port map( A => mult_143_n6022, ZN => n634);
   U521 : OAI21_X1 port map( B1 => n3675, B2 => n3645, A => n3525, ZN => 
                           mult_143_n4987);
   U522 : OAI21_X1 port map( B1 => n3675, B2 => n3596, A => mult_143_n6025, ZN 
                           => mult_143_n6024);
   U524 : OAI21_X1 port map( B1 => n3675, B2 => n3597, A => mult_143_n5889, ZN 
                           => mult_143_n5888);
   U525 : OAI21_X1 port map( B1 => n3675, B2 => n3644, A => mult_143_n5976, ZN 
                           => mult_143_n5975);
   U526 : OAI21_X1 port map( B1 => n3675, B2 => n3594, A => mult_143_n5992, ZN 
                           => mult_143_n5991);
   U530 : NOR2_X1 port map( A1 => mult_143_n6577, A2 => n2769, ZN => 
                           mult_143_n4797);
   U532 : NAND2_X1 port map( A1 => n1060, A2 => mult_143_n6118, ZN => 
                           mult_143_n6105);
   U533 : OAI21_X1 port map( B1 => mult_143_n4761, B2 => n984, A => n954, ZN =>
                           mult_143_n4759);
   U534 : OAI21_X1 port map( B1 => n1063, B2 => n984, A => n954, ZN => n817);
   U536 : OAI21_X1 port map( B1 => B_SIG(17), B2 => mult_143_n6000, A => 
                           B_SIG(18), ZN => mult_143_n6001);
   U537 : OAI21_X1 port map( B1 => B_SIG(18), B2 => n2910, A => mult_143_n6001,
                           ZN => mult_143_n5999);
   U538 : NAND2_X1 port map( A1 => B_SIG(20), A2 => n819, ZN => n818);
   U539 : OR2_X1 port map( A1 => n818, A2 => n820, ZN => mult_143_n6095);
   U540 : NOR2_X1 port map( A1 => mult_143_n6115, A2 => n826, ZN => n820);
   U541 : NOR2_X1 port map( A1 => mult_143_n5138, A2 => mult_143_n5137, ZN => 
                           n1609);
   U542 : OR2_X1 port map( A1 => mult_143_n5291, A2 => n728, ZN => n821);
   U544 : OAI21_X1 port map( B1 => mult_143_n4824, B2 => mult_143_n3007, A => 
                           mult_143_n4878, ZN => mult_143_n4877);
   U545 : OAI21_X1 port map( B1 => mult_143_n4891, B2 => mult_143_n3007, A => 
                           mult_143_n4961, ZN => mult_143_n4960);
   U546 : OAI21_X1 port map( B1 => n3645, B2 => n3656, A => mult_143_n4924, ZN 
                           => mult_143_n4923);
   U547 : OAI21_X1 port map( B1 => n3594, B2 => n3656, A => mult_143_n4861, ZN 
                           => mult_143_n4860);
   U548 : OAI21_X1 port map( B1 => mult_143_n4848, B2 => n1061, A => 
                           mult_143_n5931, ZN => mult_143_n5930);
   U550 : OAI21_X1 port map( B1 => n1061, B2 => mult_143_n5859, A => 
                           mult_143_n5880, ZN => mult_143_n5879);
   U551 : OAI21_X1 port map( B1 => n3657, B2 => n3659, A => mult_143_n5816, ZN 
                           => mult_143_n5815);
   U552 : AOI222_X1 port map( A1 => n1613, A2 => n1620, B1 => n1613, B2 => 
                           mult_143_n4869, C1 => mult_143_n4869, C2 => n1620, 
                           ZN => mult_143_n917);
   U554 : AOI222_X1 port map( A1 => n660, A2 => mult_143_n5086, B1 => 
                           mult_143_n5086, B2 => n4754, C1 => n4651, C2 => 
                           n4754, ZN => mult_143_n652);
   U559 : XNOR2_X1 port map( A => mult_143_n5309, B => n3811, ZN => 
                           mult_143_n5306);
   U562 : INV_X1 port map( A => mult_143_n5604, ZN => n699);
   U563 : AOI222_X1 port map( A1 => n3633, A2 => n3626, B1 => n3633, B2 => 
                           n3629, C1 => n3626, C2 => n3629, ZN => 
                           mult_143_n5604);
   U565 : OAI21_X1 port map( B1 => mult_143_n2458, B2 => mult_143_n4842, A => 
                           mult_143_n6295, ZN => mult_143_n6294);
   U566 : OAI222_X1 port map( A1 => n629, A2 => n978, B1 => n977, B2 => n630, 
                           C1 => mult_143_n4824, C2 => mult_143_n2458, ZN => 
                           mult_143_n6232);
   U567 : OAI222_X1 port map( A1 => n629, A2 => n979, B1 => n996, B2 => n630, 
                           C1 => mult_143_n4820, C2 => mult_143_n2458, ZN => 
                           mult_143_n6184);
   U568 : OAI222_X1 port map( A1 => n1052, A2 => n629, B1 => n981, B2 => n630, 
                           C1 => mult_143_n4828, C2 => mult_143_n2458, ZN => 
                           mult_143_n6157);
   U569 : OAI222_X1 port map( A1 => n629, A2 => n974, B1 => n976, B2 => n630, 
                           C1 => mult_143_n4848, C2 => mult_143_n2458, ZN => 
                           mult_143_n6142);
   U570 : OAI222_X1 port map( A1 => mult_143_n2458, A2 => mult_143_n5859, B1 =>
                           n1053, B2 => n630, C1 => n629, C2 => n980, ZN => 
                           mult_143_n6132);
   U571 : OAI222_X1 port map( A1 => n629, A2 => n982, B1 => n997, B2 => n630, 
                           C1 => mult_143_n4891, C2 => mult_143_n2458, ZN => 
                           mult_143_n5402);
   U572 : XNOR2_X1 port map( A => mult_143_n6232, B => A_SIG(17), ZN => 
                           mult_143_n6208);
   U573 : XNOR2_X1 port map( A => mult_143_n4844, B => mult_143_n4845, ZN => 
                           n1608);
   U574 : NOR2_X1 port map( A1 => mult_143_n4844, A2 => mult_143_n4845, ZN => 
                           mult_143_n4812);
   U576 : XNOR2_X1 port map( A => mult_143_n6208, B => mult_143_n6209, ZN => 
                           mult_143_n6204);
   U577 : NOR2_X1 port map( A1 => mult_143_n6168, A2 => mult_143_n6169, ZN => 
                           mult_143_n6173);
   U578 : XNOR2_X1 port map( A => mult_143_n6168, B => mult_143_n6169, ZN => 
                           n1607);
   U579 : NOR2_X1 port map( A1 => n1782, A2 => mult_143_n1116, ZN => 
                           mult_143_n6135);
   U580 : NOR2_X1 port map( A1 => n3695, A2 => n3526, ZN => n1606);
   U581 : AOI21_X1 port map( B1 => n3694, B2 => n3693, A => n3519, ZN => 
                           mult_143_n522);
   U582 : OAI21_X1 port map( B1 => mult_143_n4812, B2 => mult_143_n4813, A => 
                           mult_143_n4811, ZN => n1522);
   U583 : XNOR2_X1 port map( A => mult_143_n4812, B => mult_143_n4813, ZN => 
                           mult_143_n4810);
   U585 : AOI21_X1 port map( B1 => B_SIG(1), B2 => n1027, A => mult_143_n6298, 
                           ZN => mult_143_n6297);
   U586 : AOI21_X1 port map( B1 => B_SIG(1), B2 => n799, A => mult_143_n5404, 
                           ZN => mult_143_n5403);
   U587 : AOI21_X1 port map( B1 => n787, B2 => B_SIG(1), A => mult_143_n6159, 
                           ZN => mult_143_n6158);
   U588 : XNOR2_X1 port map( A => n3663, B => n3721, ZN => mult_143_n6216);
   U589 : XNOR2_X1 port map( A => mult_143_n6173, B => mult_143_n6174, ZN => 
                           mult_143_n1070);
   U590 : AOI21_X1 port map( B1 => B_SIG(1), B2 => n1023, A => mult_143_n6144, 
                           ZN => mult_143_n6143);
   U591 : OAI221_X1 port map( B1 => mult_143_n6265, B2 => A_SIG(20), C1 => 
                           mult_143_n6265, C2 => mult_143_n6266, A => 
                           mult_143_n4845, ZN => mult_143_n6261);
   U593 : AOI22_X1 port map( A1 => n3564, A2 => n3658, B1 => n4577, B2 => n4606
                           , ZN => mult_143_n6611);
   U594 : OAI222_X1 port map( A1 => n3658, A2 => n1606, B1 => n3658, B2 => 
                           n3564, C1 => n1606, C2 => n3564, ZN => 
                           mult_143_n5228);
   U595 : XNOR2_X1 port map( A => mult_143_n1536, B => mult_143_n4947, ZN => 
                           n1604);
   U601 : OAI211_X1 port map( C1 => mult_143_n6293, C2 => n629, A => A_SIG(20),
                           B => mult_143_n6265, ZN => mult_143_n4845);
   U602 : OAI21_X1 port map( B1 => n629, B2 => mult_143_n6231, A => A_SIG(17), 
                           ZN => mult_143_n6209);
   U603 : OAI21_X1 port map( B1 => n629, B2 => mult_143_n6181, A => A_SIG(14), 
                           ZN => mult_143_n6169);
   U604 : NOR2_X1 port map( A1 => n629, A2 => n643, ZN => mult_143_n1116);
   U605 : OAI21_X1 port map( B1 => n629, B2 => n641, A => A_SIG(5), ZN => 
                           mult_143_n5127);
   U606 : OAI211_X1 port map( C1 => n629, C2 => mult_143_n4832, A => n748, B =>
                           mult_143_n4831, ZN => mult_143_n4851);
   U607 : NAND4_X1 port map( A1 => A_SIG(2), A2 => n630, A3 => n910, A4 => n629
                           , ZN => mult_143_n5120);
   U608 : AOI221_X1 port map( B1 => n641, B2 => mult_143_n5120, C1 => n629, C2 
                           => mult_143_n5120, A => mult_143_n5121, ZN => 
                           mult_143_n5119);
   U609 : NOR2_X1 port map( A1 => n629, A2 => mult_143_n4832, ZN => 
                           mult_143_n4813);
   U610 : OAI21_X1 port map( B1 => n629, B2 => mult_143_n4832, A => n748, ZN =>
                           mult_143_n4830);
   U611 : NOR2_X1 port map( A1 => n629, A2 => n630, ZN => mult_143_n4555);
   U612 : OAI21_X1 port map( B1 => mult_143_n4842, B2 => mult_143_n3094, A => 
                           mult_143_n6299, ZN => mult_143_n6298);
   U613 : OAI21_X1 port map( B1 => mult_143_n4891, B2 => n2817, A => 
                           mult_143_n5405, ZN => mult_143_n5404);
   U614 : OAI21_X1 port map( B1 => mult_143_n4828, B2 => n2817, A => 
                           mult_143_n6160, ZN => mult_143_n6159);
   U615 : XNOR2_X1 port map( A => n649, B => mult_143_n6182, ZN => 
                           mult_143_n6174);
   U616 : OAI21_X1 port map( B1 => mult_143_n4848, B2 => n2817, A => 
                           mult_143_n6145, ZN => mult_143_n6144);
   U617 : XNOR2_X1 port map( A => n1612, B => A_SIG(20), ZN => mult_143_n6266);
   U618 : AOI21_X1 port map( B1 => mult_143_n6226, B2 => n3686, A => n3720, ZN 
                           => n986);
   U620 : NAND2_X1 port map( A1 => mult_143_n6146, A2 => mult_143_n6147, ZN => 
                           mult_143_n6149);
   U621 : XNOR2_X1 port map( A => mult_143_n6133, B => n642, ZN => 
                           mult_143_n5138);
   U622 : AOI21_X1 port map( B1 => n1521, B2 => n3685, A => n3748, ZN => 
                           mult_143_n1059);
   U623 : AOI21_X1 port map( B1 => mult_143_n5413, B2 => n2746, A => 
                           mult_143_n5412, ZN => mult_143_n1101);
   U625 : AOI22_X1 port map( A1 => mult_143_n1863, A2 => n686, B1 => 
                           mult_143_n1123, B2 => n693, ZN => mult_143_n4947);
   U631 : OAI21_X1 port map( B1 => mult_143_n6029, B2 => n1072, A => 
                           mult_143_n5940, ZN => mult_143_n6129);
   U634 : AOI22_X1 port map( A1 => n3827, A2 => n3820, B1 => n3779, B2 => n3772
                           , ZN => mult_143_n5009);
   U635 : AOI22_X1 port map( A1 => B_SIG(4), A2 => mult_143_n96, B1 => B_SIG(6)
                           , B2 => n2598, ZN => mult_143_n4892);
   U636 : AOI22_X1 port map( A1 => n3782, A2 => n3820, B1 => n3783, B2 => n3772
                           , ZN => mult_143_n5047);
   U638 : AOI22_X1 port map( A1 => n3779, A2 => n3531, B1 => n3781, B2 => n4677
                           , ZN => mult_143_n5018);
   U640 : AOI22_X1 port map( A1 => n3787, A2 => n3531, B1 => n3789, B2 => n3772
                           , ZN => mult_143_n6101);
   U641 : AOI22_X1 port map( A1 => n4871, A2 => n3531, B1 => n4765, B2 => n3772
                           , ZN => mult_143_n6109);
   U642 : OAI21_X1 port map( B1 => n3664, B2 => n3643, A => mult_143_n5009, ZN 
                           => mult_143_n5008);
   U660 : AOI22_X1 port map( A1 => B_SIG(4), A2 => n772, B1 => B_SIG(2), B2 => 
                           mult_143_n72, ZN => mult_143_n6275);
   U661 : AOI22_X1 port map( A1 => B_SIG(3), A2 => mult_143_n3245, B1 => 
                           B_SIG(2), B2 => n1030, ZN => mult_143_n5131);
   U662 : AOI22_X1 port map( A1 => B_SIG(4), A2 => n765, B1 => B_SIG(2), B2 => 
                           mult_143_n48, ZN => mult_143_n6172);
   U663 : AOI22_X1 port map( A1 => B_SIG(4), A2 => n2599, B1 => B_SIG(2), B2 =>
                           mult_143_n6621, ZN => mult_143_n6207);
   U664 : AOI22_X1 port map( A1 => B_SIG(1), A2 => mult_143_n36, B1 => B_SIG(2)
                           , B2 => n1023, ZN => mult_143_n6141);
   U668 : AOI21_X1 port map( B1 => B_SIG(5), B2 => n799, A => mult_143_n4890, 
                           ZN => mult_143_n4889);
   U669 : OAI21_X1 port map( B1 => B_SIG(5), B2 => B_SIG(3), A => B_SIG(4), ZN 
                           => mult_143_n6288);
   U671 : NAND2_X1 port map( A1 => mult_143_n6105, A2 => mult_143_n6106, ZN => 
                           mult_143_n6102);
   U673 : XNOR2_X1 port map( A => mult_143_n6102, B => mult_143_n6103, ZN => 
                           mult_143_n4407);
   U675 : XOR2_X1 port map( A => mult_143_n6026, B => B_SIG(15), Z => 
                           mult_143_n2981);
   U677 : OAI21_X1 port map( B1 => mult_143_n4842, B2 => mult_143_n6624, A => 
                           mult_143_n5028, ZN => mult_143_n5027);
   U678 : OAI21_X1 port map( B1 => mult_143_n4824, B2 => n1075, A => 
                           mult_143_n4971, ZN => mult_143_n4970);
   U679 : OAI21_X1 port map( B1 => n3673, B2 => n3653, A => mult_143_n4858, ZN 
                           => mult_143_n4857);
   U680 : OAI21_X1 port map( B1 => n3644, B2 => n3652, A => mult_143_n4875, ZN 
                           => mult_143_n4874);
   U681 : OAI21_X1 port map( B1 => n3643, B2 => n3653, A => mult_143_n6083, ZN 
                           => mult_143_n6082);
   U682 : OAI21_X1 port map( B1 => n3594, B2 => n3652, A => mult_143_n5995, ZN 
                           => mult_143_n5994);
   U683 : OAI21_X1 port map( B1 => n3653, B2 => n3597, A => mult_143_n5895, ZN 
                           => mult_143_n5894);
   U684 : OAI21_X1 port map( B1 => n1075, B2 => mult_143_n5124, A => 
                           mult_143_n5834, ZN => mult_143_n5833);
   U685 : OAI221_X1 port map( B1 => mult_143_n6122, B2 => mult_143_n6106, C1 =>
                           mult_143_n6122, C2 => mult_143_n6105, A => 
                           mult_143_n6123, ZN => mult_143_n6120);
   U688 : AOI22_X1 port map( A1 => n3646, A2 => n3766, B1 => n3540, B2 => n3827
                           , ZN => mult_143_n4954);
   U689 : AOI22_X1 port map( A1 => n778, A2 => B_SIG(15), B1 => mult_143_n84, 
                           B2 => B_SIG(13), ZN => mult_143_n4988);
   U690 : AOI21_X1 port map( B1 => n3819, B2 => n3800, A => mult_143_n4926, ZN 
                           => mult_143_n4925);
   U692 : AOI22_X1 port map( A1 => B_SIG(4), A2 => mult_143_n48, B1 => B_SIG(6)
                           , B2 => n765, ZN => mult_143_n6191);
   U693 : AOI22_X1 port map( A1 => B_SIG(4), A2 => mult_143_n72, B1 => B_SIG(6)
                           , B2 => n772, ZN => mult_143_n4825);
   U694 : AOI22_X1 port map( A1 => B_SIG(4), A2 => mult_143_n6621, B1 => 
                           B_SIG(6), B2 => n2599, ZN => mult_143_n6248);
   U695 : AOI22_X1 port map( A1 => B_SIG(4), A2 => mult_143_n36, B1 => B_SIG(6)
                           , B2 => n755, ZN => mult_143_n5922);
   U696 : AOI21_X1 port map( B1 => B_SIG(4), B2 => n2598, A => mult_143_n6069, 
                           ZN => mult_143_n6068);
   U697 : AOI21_X1 port map( B1 => B_SIG(4), B2 => n799, A => mult_143_n6072, 
                           ZN => mult_143_n6071);
   U703 : AOI21_X1 port map( B1 => n3800, B2 => n3807, A => mult_143_n4863, ZN 
                           => mult_143_n4862);
   U704 : AOI21_X1 port map( B1 => n3800, B2 => n4665, A => mult_143_n4880, ZN 
                           => mult_143_n4879);
   U705 : AOI22_X1 port map( A1 => B_SIG(11), A2 => mult_143_n72, B1 => 
                           B_SIG(13), B2 => n772, ZN => mult_143_n6020);
   U706 : AOI21_X1 port map( B1 => B_SIG(13), B2 => n1027, A => mult_143_n4963,
                           ZN => mult_143_n4962);
   U708 : AOI22_X1 port map( A1 => B_SIG(11), A2 => mult_143_n3228, B1 => 
                           B_SIG(13), B2 => n1026, ZN => mult_143_n5883);
   U709 : AOI22_X1 port map( A1 => n3827, A2 => n3799, B1 => n3800, B2 => n3823
                           , ZN => mult_143_n5934);
   U710 : AOI21_X1 port map( B1 => n3780, B2 => n3802, A => mult_143_n5972, ZN 
                           => mult_143_n5971);
   U711 : AOI21_X1 port map( B1 => n778, B2 => B_SIG(3), A => mult_143_n4841, 
                           ZN => mult_143_n4840);
   U712 : AOI21_X1 port map( B1 => n774, B2 => B_SIG(3), A => mult_143_n6274, 
                           ZN => mult_143_n6273);
   U713 : AOI21_X1 port map( B1 => n787, B2 => B_SIG(3), A => mult_143_n6171, 
                           ZN => mult_143_n6170);
   U714 : AOI21_X1 port map( B1 => n765, B2 => B_SIG(3), A => mult_143_n6155, 
                           ZN => mult_143_n6154);
   U715 : AOI22_X1 port map( A1 => n778, A2 => B_SIG(5), B1 => mult_143_n84, B2
                           => B_SIG(3), ZN => mult_143_n6053);
   U716 : AOI22_X1 port map( A1 => n1027, A2 => B_SIG(3), B1 => mult_143_n84, 
                           B2 => B_SIG(2), ZN => mult_143_n6050);
   U718 : NAND2_X1 port map( A1 => mult_143_n5291, A2 => n728, ZN => 
                           mult_143_n5296);
   U722 : AND2_X1 port map( A1 => n813, A2 => n814, ZN => n943);
   U738 : INV_X1 port map( A => mult_143_n5250, ZN => n702);
   U741 : INV_X1 port map( A => mult_143_n5747, ZN => n717);
   U742 : INV_X1 port map( A => mult_143_n5470, ZN => n718);
   U743 : INV_X1 port map( A => mult_143_n5418, ZN => n714);
   U745 : INV_X1 port map( A => mult_143_n5586, ZN => n730);
   U746 : INV_X1 port map( A => mult_143_n5677, ZN => n734);
   U749 : AOI222_X1 port map( A1 => n4864, A2 => n4758, B1 => n3104, B2 => 
                           mult_143_n5401, C1 => n4758, C2 => mult_143_n5401, 
                           ZN => n1480);
   U752 : AOI221_X1 port map( B1 => B_SIG(5), B2 => n1031, C1 => B_SIG(4), C2 
                           => mult_143_n3228, A => mult_143_n5865, ZN => 
                           mult_143_n5864);
   U759 : INV_X1 port map( A => mult_143_n4774, ZN => n747);
   U760 : INV_X1 port map( A => mult_143_n4777, ZN => n727);
   U761 : INV_X1 port map( A => mult_143_n4775, ZN => n726);
   U768 : INV_X1 port map( A => mult_143_n6029, ZN => n636);
   U778 : INV_X1 port map( A => mult_143_n4788, ZN => n721);
   U789 : OR2_X1 port map( A1 => mult_143_n6199, A2 => mult_143_n6200, ZN => 
                           n980);
   U792 : AND4_X1 port map( A1 => n4936, A2 => mult_143_n4401, A3 => n2936, A4 
                           => n4901, ZN => n824);
   U803 : INV_X1 port map( A => mult_143_n5787, ZN => n712);
   U805 : INV_X1 port map( A => mult_143_n1528, ZN => n667);
   U806 : INV_X1 port map( A => mult_143_n6293, ZN => n651);
   U816 : INV_X1 port map( A => mult_143_n1537, ZN => n1832);
   U831 : OR2_X1 port map( A1 => mult_143_n6148, A2 => mult_143_n6149, ZN => 
                           n1601);
   U832 : INV_X1 port map( A => mult_143_n6181, ZN => n648);
   U839 : INV_X1 port map( A => n2824, ZN => n631);
   U845 : XOR2_X1 port map( A => mult_143_n6285, B => n825, Z => mult_143_n2919
                           );
   U851 : INV_X1 port map( A => mult_143_n5316, ZN => n728);
   U856 : INV_X1 port map( A => mult_143_n6231, ZN => n650);
   U858 : OR2_X1 port map( A1 => mult_143_n6306, A2 => mult_143_n6231, ZN => 
                           n977);
   U859 : INV_X1 port map( A => n977, ZN => n772);
   U865 : OR2_X1 port map( A1 => mult_143_n6284, A2 => mult_143_n6181, ZN => 
                           n996);
   U871 : OR2_X1 port map( A1 => n3721, A2 => n3663, ZN => mult_143_n6226);
   U885 : INV_X1 port map( A => mult_143_n6254, ZN => n643);
   U889 : OR2_X1 port map( A1 => mult_143_n6253, A2 => n643, ZN => n976);
   U895 : INV_X1 port map( A => mult_143_n6199, ZN => n641);
   U903 : INV_X1 port map( A => A_SIG(1), ZN => n639);
   U904 : INV_X1 port map( A => A_SIG(0), ZN => n638);
   U930 : OR3_X1 port map( A1 => n3715, A2 => n3677, A3 => n3558, ZN => n1521);
   U931 : INV_X1 port map( A => mult_143_n6098, ZN => n819);
   U932 : AND2_X1 port map( A1 => n3787, A2 => n3807, ZN => n811);
   U937 : OR2_X1 port map( A1 => mult_143_n5128, A2 => mult_143_n5127, ZN => 
                           mult_143_n5137);
   U946 : INV_X1 port map( A => mult_143_n1818, ZN => n1828);
   U950 : INV_X1 port map( A => n976, ZN => n755);
   U954 : INV_X1 port map( A => mult_143_n1123, ZN => n686);
   U955 : INV_X1 port map( A => mult_143_n1863, ZN => n693);
   U960 : INV_X1 port map( A => mult_143_n1815, ZN => n688);
   U962 : INV_X1 port map( A => mult_143_n5084, ZN => n680);
   U968 : NAND2_X1 port map( A1 => mult_143_n5303, A2 => mult_143_n5304, ZN => 
                           n1003);
   U970 : NAND2_X1 port map( A1 => n1003, A2 => n2736, ZN => n1005);
   U971 : OAI211_X1 port map( C1 => mult_143_n5303, C2 => mult_143_n5304, A => 
                           n1005, B => mult_143_n5305, ZN => mult_143_n5299);
   U977 : NAND2_X1 port map( A1 => mult_143_n5306, A2 => n3640, ZN => n1010);
   U981 : NAND2_X1 port map( A1 => n1010, A2 => n1013, ZN => mult_143_n5307);
   U986 : INV_X1 port map( A => mw_I4sum_7_port, ZN => EXP_in(7));
   U109 : NOR2_X1 port map( A1 => mult_143_n5040, A2 => n431, ZN => n1600);
   U101 : INV_X1 port map( A => B_SIG(17), ZN => n423);
   mult_143_U4012 : XNOR2_X1 port map( A => A_SIG(18), B => A_SIG(19), ZN => 
                           mult_143_n6301);
   mult_143_U4022 : XNOR2_X1 port map( A => A_SIG(16), B => A_SIG(15), ZN => 
                           mult_143_n6305);
   mult_143_U3935 : XNOR2_X1 port map( A => A_SIG(9), B => A_SIG(10), ZN => 
                           mult_143_n6242);
   mult_143_U3996 : XNOR2_X1 port map( A => A_SIG(12), B => A_SIG(13), ZN => 
                           mult_143_n6292);
   mult_143_U3960 : XNOR2_X1 port map( A => A_SIG(7), B => A_SIG(6), ZN => 
                           mult_143_n6255);
   mult_143_U4675 : XOR2_X1 port map( A => A_SIG(15), B => n649, Z => 
                           mult_143_n6231);
   U797 : OR2_X1 port map( A1 => mult_143_n6254, A2 => mult_143_n6255, ZN => 
                           n974);
   mult_143_U4668 : XOR2_X1 port map( A => n1765, B => A_SIG(12), Z => 
                           mult_143_n6181);
   U400 : INV_X1 port map( A => mult_143_n4832, ZN => n654);
   U887 : NAND2_X1 port map( A1 => mult_143_n6254, A2 => mult_143_n6253, ZN => 
                           mult_143_n4848);
   U197 : NAND2_X1 port map( A1 => n886, A2 => B_SIG(7), ZN => n487);
   U484 : OR2_X1 port map( A1 => n895, A2 => n891, ZN => n808);
   U366 : NAND2_X1 port map( A1 => n2778, A2 => n2634, ZN => n603);
   mult_143_U2420 : NAND2_X1 port map( A1 => n2855, A2 => n2603, ZN => 
                           mult_143_n4768);
   mult_143_U2883 : NOR2_X1 port map( A1 => n1725, A2 => n1755, ZN => 
                           mult_143_n5312);
   mult_143_U2884 : AOI21_X1 port map( B1 => n1755, B2 => n1725, A => n1743, ZN
                           => mult_143_n5311);
   mult_143_U2886 : XNOR2_X1 port map( A => n3617, B => n3623, ZN => 
                           mult_143_n5313);
   U295 : XNOR2_X1 port map( A => n4611, B => n4608, ZN => n555);
   U88 : NAND2_X1 port map( A1 => n2696, A2 => n3065, ZN => n415);
   mult_143_U3217 : AOI222_X1 port map( A1 => n2727, A2 => n2669, B1 => n2727, 
                           B2 => n2691, C1 => n2669, C2 => n2691, ZN => 
                           mult_143_n5174);
   U212 : NAND2_X1 port map( A1 => n2695, A2 => mult_143_n6572, ZN => n496);
   mult_143_U3185 : AOI222_X1 port map( A1 => n3630, A2 => n4633, B1 => n3630, 
                           B2 => n3619, C1 => n4633, C2 => n3619, ZN => 
                           mult_143_n5631);
   U978 : NAND2_X1 port map( A1 => n3618, A2 => n1718, ZN => n1011);
   mult_143_U2901 : XNOR2_X1 port map( A => n3638, B => n3764, ZN => 
                           mult_143_n5326);
   mult_143_U2913 : XNOR2_X1 port map( A => n3637, B => n3635, ZN => 
                           mult_143_n5337);
   mult_143_U2911 : AOI21_X1 port map( B1 => n3638, B2 => n3764, A => n3624, ZN
                           => mult_143_n5335);
   U271 : NOR2_X1 port map( A1 => B_SIG(9), A2 => n878, ZN => n538);
   U836 : XOR2_X1 port map( A => A_SIG(23), B => A_SIG(22), Z => mult_143_n6110
                           );
   U833 : OR2_X1 port map( A1 => n654, A2 => mult_143_n6111, ZN => n982);
   U980 : NAND2_X1 port map( A1 => n1011, A2 => n3761, ZN => n1013);
   mult_143_U2900 : XNOR2_X1 port map( A => mult_143_n5326, B => n3624, ZN => 
                           mult_143_n5321);
   mult_143_U2912 : XNOR2_X1 port map( A => mult_143_n5337, B => n1758, ZN => 
                           mult_143_n5330);
   mult_143_U2909 : NOR2_X1 port map( A1 => mult_143_n5335, A2 => 
                           mult_143_n5336, ZN => mult_143_n5331);
   mult_143_U2921 : XNOR2_X1 port map( A => mult_143_n5342, B => n4587, ZN => 
                           mult_143_n5334);
   mult_143_U2917 : XNOR2_X1 port map( A => mult_143_n5340, B => n3621, ZN => 
                           mult_143_n5275);
   U408 : INV_X1 port map( A => mult_143_n5341, ZN => n715);
   mult_143_U2885 : XNOR2_X1 port map( A => mult_143_n5313, B => n3639, ZN => 
                           mult_143_n5297);
   mult_143_U2882 : NOR2_X1 port map( A1 => mult_143_n5311, A2 => 
                           mult_143_n5312, ZN => mult_143_n5298);
   U119 : XNOR2_X1 port map( A => mult_143_n5315, B => n438, ZN => 
                           mult_143_n5293);
   mult_143_U3169 : XNOR2_X1 port map( A => n3814, B => mult_143_n5622, ZN => 
                           mult_143_n5601);
   U86 : NAND2_X1 port map( A1 => n415, A2 => n4632, ZN => n413);
   mult_143_U3313 : XNOR2_X1 port map( A => n3803, B => mult_143_n5746, ZN => 
                           mult_143_n5720);
   U93 : INV_X1 port map( A => mult_143_n5631, ZN => n711);
   U308 : NOR2_X1 port map( A1 => mult_143_n5735, A2 => mult_143_n5736, ZN => 
                           mult_143_n5705);
   U364 : NAND2_X1 port map( A1 => n603, A2 => n1039, ZN => n601);
   U723 : OR2_X1 port map( A1 => n650, A2 => mult_143_n6305, ZN => n978);
   U876 : INV_X1 port map( A => n982, ZN => n799);
   U837 : OR2_X1 port map( A1 => mult_143_n6110, A2 => mult_143_n4832, ZN => 
                           n997);
   mult_143_U2871 : NAND2_X1 port map( A1 => mult_143_n5293, A2 => 
                           mult_143_n5294, ZN => mult_143_n5300);
   mult_143_U2873 : NAND2_X1 port map( A1 => mult_143_n5297, A2 => n3672, ZN =>
                           mult_143_n5305);
   U223 : INV_X1 port map( A => mult_143_n5333, ZN => n506);
   mult_143_U2899 : AOI222_X1 port map( A1 => n3726, A2 => n1749, B1 => n3726, 
                           B2 => mult_143_n5321, C1 => n1749, C2 => 
                           mult_143_n5321, ZN => mult_143_n5289);
   mult_143_U2907 : XNOR2_X1 port map( A => mult_143_n5334, B => n2725, ZN => 
                           mult_143_n5332);
   mult_143_U2908 : AOI222_X1 port map( A1 => n2612, A2 => mult_143_n5330, B1 
                           => n2612, B2 => mult_143_n5331, C1 => mult_143_n5330
                           , C2 => mult_143_n5331, ZN => mult_143_n5325);
   U163 : AND2_X1 port map( A1 => mult_143_n5720, A2 => mult_143_n5719, ZN => 
                           n465);
   mult_143_U2905 : XNOR2_X1 port map( A => mult_143_n5330, B => mult_143_n5331
                           , ZN => mult_143_n5329);
   mult_143_U3333 : AOI222_X1 port map( A1 => mult_143_n5741, A2 => 
                           mult_143_n5742, B1 => mult_143_n5741, B2 => 
                           mult_143_n5743, C1 => mult_143_n5743, C2 => 
                           mult_143_n5742, ZN => mult_143_n5467);
   U363 : OAI21_X1 port map( B1 => n2778, B2 => n2634, A => n601, ZN => 
                           mult_143_n5662);
   U248 : INV_X1 port map( A => mult_143_n5297, ZN => n525);
   U294 : XNOR2_X1 port map( A => mult_143_n5290, B => n555, ZN => 
                           mult_143_n5291);
   U85 : OAI21_X1 port map( B1 => n3065, B2 => n2696, A => n413, ZN => 
                           mult_143_n5758);
   U252 : AND2_X1 port map( A1 => n3805, A2 => n3787, ZN => n528);
   U195 : NAND2_X1 port map( A1 => mult_143_n72, A2 => B_SIG(7), ZN => n486);
   U183 : AND2_X1 port map( A1 => n3539, A2 => n3787, ZN => n478);
   U209 : AND2_X1 port map( A1 => n3531, A2 => n3800, ZN => n494);
   U892 : INV_X1 port map( A => n978, ZN => n774);
   U358 : NAND2_X1 port map( A1 => n3539, A2 => n4714, ZN => n595);
   U246 : NAND2_X1 port map( A1 => n525, A2 => n4594, ZN => n523);
   U239 : NAND2_X1 port map( A1 => mult_143_n5465, A2 => mult_143_n5466, ZN => 
                           n515);
   mult_143_U2852 : AOI222_X1 port map( A1 => n1046, A2 => mult_143_n5253, B1 
                           => n1046, B2 => mult_143_n5254, C1 => mult_143_n5253
                           , C2 => mult_143_n5254, ZN => n1479);
   U94 : NAND2_X1 port map( A1 => n421, A2 => n418, ZN => mult_143_n5596);
   U222 : XNOR2_X1 port map( A => mult_143_n5332, B => n506, ZN => 
                           mult_143_n5324);
   U162 : OAI22_X1 port map( A1 => mult_143_n5718, A2 => n465, B1 => 
                           mult_143_n5720, B2 => mult_143_n5719, ZN => 
                           mult_143_n5732);
   U156 : AND2_X1 port map( A1 => n3772, A2 => n4688, ZN => n461);
   U115 : NOR2_X1 port map( A1 => n533, A2 => n435, ZN => n434);
   U76 : NAND2_X1 port map( A1 => mult_143_n5094, A2 => n408, ZN => n407);
   U110 : AND2_X1 port map( A1 => n3819, A2 => n3787, ZN => n431);
   mult_143_U3328 : AOI222_X1 port map( A1 => n698, A2 => n4950, B1 => n698, B2
                           => n2664, C1 => n2664, C2 => n3048, ZN => 
                           mult_143_n5513);
   U387 : XNOR2_X1 port map( A => mult_143_n5588, B => mult_143_n5587, ZN => 
                           n617);
   mult_143_U3259 : XNOR2_X1 port map( A => mult_143_n5694, B => mult_143_n5693
                           , ZN => mult_143_n5680);
   mult_143_U2898 : NAND2_X1 port map( A1 => mult_143_n5288, A2 => 
                           mult_143_n5289, ZN => mult_143_n5278);
   mult_143_U2896 : AOI22_X1 port map( A1 => mult_143_n5322, A2 => n4732, B1 =>
                           mult_143_n5324, B2 => mult_143_n5325, ZN => 
                           mult_143_n5280);
   mult_143_U2856 : OAI22_X1 port map( A1 => n2881, A2 => mult_143_n5261, B1 =>
                           mult_143_n5263, B2 => mult_143_n5264, ZN => 
                           mult_143_n5259);
   U342 : NOR2_X1 port map( A1 => n4955, A2 => mult_143_n5278, ZN => n583);
   U236 : NAND2_X1 port map( A1 => n514, A2 => n513, ZN => n1596);
   U159 : OAI21_X1 port map( B1 => n716, B2 => n464, A => n463, ZN => n1517);
   U47 : AOI21_X1 port map( B1 => mult_143_n5262, B2 => mult_143_n5261, A => 
                           n386, ZN => mult_143_n5267);
   U428 : XOR2_X1 port map( A => n882, B => mult_143_n6245, Z => mult_143_n6628
                           );
   U268 : INV_X1 port map( A => mult_143_n5970, ZN => n633);
   mult_143_U2467 : XNOR2_X1 port map( A => A_SIG(20), B => mult_143_n4840, ZN 
                           => mult_143_n4811);
   U270 : NAND2_X1 port map( A1 => mult_143_n5970, A2 => n538, ZN => n537);
   U411 : INV_X1 port map( A => mult_143_n5733, ZN => n1787);
   mult_143_U3024 : XNOR2_X1 port map( A => n3711, B => n3670, ZN => 
                           mult_143_n5456);
   mult_143_U2854 : NAND2_X1 port map( A1 => mult_143_n5259, A2 => 
                           mult_143_n5260, ZN => mult_143_n5258);
   mult_143_U2926 : OAI21_X1 port map( B1 => mult_143_n5265, B2 => 
                           mult_143_n5266, A => mult_143_n5267, ZN => 
                           mult_143_n5255);
   mult_143_U2969 : NAND2_X1 port map( A1 => n3595, A2 => n3606, ZN => n1594);
   U340 : NOR2_X1 port map( A1 => n583, A2 => n582, ZN => n581);
   U173 : AOI22_X1 port map( A1 => n633, A2 => B_SIG(9), B1 => n882, B2 => 
                           mult_143_n5970, ZN => n471);
   mult_143_U3201 : NOR2_X1 port map( A1 => mult_143_n5641, A2 => n4710, ZN => 
                           mult_143_n5640);
   U64 : NAND2_X1 port map( A1 => n634, A2 => n398, ZN => n397);
   U205 : XNOR2_X1 port map( A => n3095, B => mult_143_n5938, ZN => 
                           mult_143_n3443);
   U171 : XNOR2_X1 port map( A => n471, B => B_SIG(10), ZN => mult_143_n6627);
   U292 : XNOR2_X1 port map( A => n3712, B => n4621, ZN => n553);
   mult_143_U2986 : NOR2_X1 port map( A1 => n2911, A2 => mult_143_n5209, ZN => 
                           mult_143_n2868);
   mult_143_U3262 : NAND2_X1 port map( A1 => mult_143_n5696, A2 => 
                           mult_143_n5697, ZN => mult_143_n5205);
   mult_143_U3263 : NOR2_X1 port map( A1 => mult_143_n5696, A2 => 
                           mult_143_n5697, ZN => mult_143_n5204);
   U17 : INV_X1 port map( A => mult_143_n5240, ZN => n505);
   mult_143_U2793 : NAND2_X1 port map( A1 => mult_143_n5169, A2 => 
                           mult_143_n5168, ZN => mult_143_n373);
   U63 : OAI21_X1 port map( B1 => n634, B2 => n400, A => n397, ZN => n396);
   U122 : XNOR2_X1 port map( A => n440, B => mult_143_n6089, ZN => 
                           mult_143_n3137);
   mult_143_U2464 : OAI21_X1 port map( B1 => mult_143_n6627, B2 => 
                           mult_143_n4820, A => mult_143_n4839, ZN => 
                           mult_143_n4838);
   mult_143_U2824 : OAI21_X1 port map( B1 => n4882, B2 => mult_143_n344, A => 
                           mult_143_n5205, ZN => mult_143_n335);
   mult_143_U2778 : NAND2_X1 port map( A1 => mult_143_n3154, A2 => n4887, ZN =>
                           mult_143_n392);
   U62 : XNOR2_X1 port map( A => n396, B => B_SIG(13), ZN => mult_143_n3010);
   mult_143_U2463 : AOI21_X1 port map( B1 => B_SIG(10), B2 => n2599, A => 
                           mult_143_n4838, ZN => mult_143_n4837);
   mult_143_U2482 : AOI21_X1 port map( B1 => n3778, B2 => n4665, A => 
                           mult_143_n4860, ZN => mult_143_n4859);
   U368 : OAI21_X1 port map( B1 => n605, B2 => mult_143_n4502, A => n604, ZN =>
                           mult_143_n3055);
   U45 : XNOR2_X1 port map( A => n3544, B => n3812, ZN => SIG_in(27));
   mult_143_U2481 : XNOR2_X1 port map( A => mult_143_n4859, B => n3773, ZN => 
                           n1590);
   mult_143_U2560 : AOI21_X1 port map( B1 => n4695, B2 => n3805, A => n3542, ZN
                           => mult_143_n4941);
   mult_143_U2810 : AOI21_X1 port map( B1 => B_SIG(14), B2 => mult_143_n6621, A
                           => mult_143_n5193, ZN => mult_143_n5192);
   U315 : AOI21_X1 port map( B1 => n567, B2 => n566, A => n564, ZN => 
                           mult_143_n4846);
   mult_143_U2821 : OAI21_X1 port map( B1 => n3644, B2 => n1584, A => 
                           mult_143_n5203, ZN => mult_143_n5201);
   mult_143_U3043 : AOI222_X1 port map( A1 => n1677, A2 => n3698, B1 => n1677, 
                           B2 => n3697, C1 => n3698, C2 => n3697, ZN => 
                           mult_143_n2702);
   mult_143_U3609 : OAI21_X1 port map( B1 => n3594, B2 => n1589, A => 
                           mult_143_n2133, ZN => mult_143_n6008);
   mult_143_U3713 : OAI21_X1 port map( B1 => n1584, B2 => n3645, A => n3055, ZN
                           => mult_143_n6066);
   mult_143_U3681 : OAI21_X1 port map( B1 => n3596, B2 => n1589, A => 
                           mult_143_n2066, ZN => mult_143_n6047);
   mult_143_U3781 : OAI21_X1 port map( B1 => n1584, B2 => n3643, A => n3068, ZN
                           => mult_143_n6119);
   mult_143_U2625 : AOI21_X1 port map( B1 => B_SIG(11), B2 => mult_143_n96, A 
                           => mult_143_n5001, ZN => n1515);
   mult_143_U3558 : OAI21_X1 port map( B1 => n3673, B2 => n1589, A => 
                           mult_143_n2267, ZN => mult_143_n5960);
   mult_143_U3510 : OAI21_X1 port map( B1 => n3597, B2 => n1584, A => n3063, ZN
                           => mult_143_n5914);
   mult_143_U2809 : XNOR2_X1 port map( A => n3773, B => n3552, ZN => n1588);
   U82 : XNOR2_X1 port map( A => n3546, B => n2780, ZN => mult_143_n5050);
   mult_143_U2614 : XNOR2_X1 port map( A => mult_143_n4991, B => n2864, ZN => 
                           mult_143_n4989);
   mult_143_U2576 : XNOR2_X1 port map( A => mult_143_n4957, B => mult_143_n4956
                           , ZN => n970);
   U155 : NOR2_X1 port map( A1 => mult_143_n5080, A2 => n461, ZN => n460);
   U132 : NOR2_X1 port map( A1 => mult_143_n5948, A2 => n446, ZN => n445);
   U189 : AND2_X1 port map( A1 => n1572, A2 => n4630, ZN => n482);
   mult_143_U2820 : XNOR2_X1 port map( A => mult_143_n5201, B => n4754, ZN => 
                           n955);
   U182 : NOR2_X1 port map( A1 => mult_143_n5199, A2 => n478, ZN => n1587);
   U154 : XNOR2_X1 port map( A => n460, B => n4752, ZN => mult_143_n5075);
   U180 : XNOR2_X1 port map( A => n1587, B => n3795, ZN => mult_143_n3455);
   mult_143_U3435 : AOI21_X1 port map( B1 => n3789, B2 => n3801, A => n1523, ZN
                           => mult_143_n5847);
   mult_143_U3551 : AOI21_X1 port map( B1 => n4714, B2 => n3817, A => n3560, ZN
                           => mult_143_n5953);
   U924 : INV_X1 port map( A => B_SIG(20), ZN => n851);
   mult_143_U2893 : XNOR2_X1 port map( A => n3688, B => n3620, ZN => 
                           mult_143_n5290);
   U262 : AND2_X1 port map( A1 => n3806, A2 => n3786, ZN => n533);
   U639 : AOI221_X1 port map( B1 => n2598, B2 => B_SIG(3), C1 => B_SIG(1), C2 
                           => mult_143_n96, A => mult_143_n5231, ZN => 
                           mult_143_n5230);
   U49 : XNOR2_X1 port map( A => n387, B => n1046, ZN => mult_143_n5262);
   mult_143_U2506 : AOI21_X1 port map( B1 => B_SIG(8), B2 => n1027, A => 
                           mult_143_n4887, ZN => mult_143_n4886);
   U75 : AOI21_X1 port map( B1 => n3641, B2 => n4672, A => n407, ZN => 
                           mult_143_n5092);
   mult_143_U3803 : AOI21_X1 port map( B1 => B_SIG(19), B2 => B_SIG(17), A => 
                           B_SIG(18), ZN => mult_143_n6115);
   mult_143_U2866 : AOI222_X1 port map( A1 => n4611, A2 => n4608, B1 => n4611, 
                           B2 => mult_143_n5290, C1 => n4608, C2 => 
                           mult_143_n5290, ZN => mult_143_n5285);
   U334 : AOI222_X1 port map( A1 => n4618, A2 => n4613, B1 => n4618, B2 => 
                           n3811, C1 => n4613, C2 => n3811, ZN => 
                           mult_143_n5304);
   mult_143_U2860 : AOI222_X1 port map( A1 => n715, A2 => mult_143_n5275, B1 =>
                           n715, B2 => mult_143_n5276, C1 => mult_143_n5275, C2
                           => mult_143_n5276, ZN => mult_143_n5269);
   U253 : AND2_X1 port map( A1 => mult_143_n5296, A2 => n545, ZN => n544);
   U7 : AND2_X1 port map( A1 => B_SIG(5), A2 => B_SIG(7), ZN => n1018);
   U11 : NAND2_X1 port map( A1 => mult_143_n6272, A2 => n1018, ZN => n1070);
   U12 : OAI21_X1 port map( B1 => n2895, B2 => n4651, A => n1019, ZN => 
                           mult_143_n5087);
   U14 : NAND2_X1 port map( A1 => n660, A2 => n2895, ZN => n1019);
   U22 : INV_X1 port map( A => n974, ZN => n1023);
   U26 : AOI222_X1 port map( A1 => n3650, A2 => n3711, B1 => n3650, B2 => n3670
                           , C1 => n3711, C2 => n3670, ZN => mult_143_n5434);
   U27 : AOI222_X1 port map( A1 => mult_143_n5424, A2 => mult_143_n5425, B1 => 
                           mult_143_n5424, B2 => n724, C1 => n724, C2 => 
                           mult_143_n5425, ZN => n1477);
   U33 : AOI222_X1 port map( A1 => mult_143_n5725, A2 => n4858, B1 => 
                           mult_143_n5725, B2 => mult_143_n5728, C1 => n4858, 
                           C2 => mult_143_n5728, ZN => mult_143_n5469);
   U34 : AOI222_X1 port map( A1 => n699, A2 => mult_143_n4361, B1 => n699, B2 
                           => n2609, C1 => mult_143_n4361, C2 => n2609, ZN => 
                           n1066);
   U57 : XNOR2_X1 port map( A => n634, B => mult_143_n6256, ZN => 
                           mult_143_n6626);
   U58 : OR2_X1 port map( A1 => mult_143_n6208, A2 => mult_143_n6209, ZN => 
                           n1579);
   U66 : AOI222_X1 port map( A1 => n4729, A2 => mult_143_n5514, B1 => 
                           mult_143_n5513, B2 => mult_143_n5515, C1 => 
                           mult_143_n5514, C2 => mult_143_n5515, ZN => n1475);
   U68 : XOR2_X1 port map( A => n632, B => mult_143_n6249, Z => mult_143_n2800)
                           ;
   U70 : OR2_X1 port map( A1 => mult_143_n5722, A2 => mult_143_n5723, ZN => 
                           n562);
   U105 : INV_X1 port map( A => mult_143_n6115, ZN => n1032);
   U108 : XNOR2_X1 port map( A => n1755, B => n1725, ZN => mult_143_n5310);
   U112 : XNOR2_X1 port map( A => n1651, B => n3615, ZN => n438);
   U117 : OR2_X1 port map( A1 => mult_143_n5293, A2 => mult_143_n5294, ZN => 
                           n545);
   U118 : NOR2_X1 port map( A1 => n3764, A2 => n3638, ZN => mult_143_n5336);
   U120 : NOR2_X1 port map( A1 => mult_143_n5322, A2 => n4732, ZN => 
                           mult_143_n5279);
   U121 : NOR2_X1 port map( A1 => mult_143_n5280, A2 => mult_143_n5279, ZN => 
                           n582);
   U129 : AOI222_X1 port map( A1 => mult_143_n6435, A2 => n1752, B1 => 
                           mult_143_n6435, B2 => n1731, C1 => n1752, C2 => 
                           n1731, ZN => mult_143_n5352);
   U130 : AND2_X1 port map( A1 => mult_143_n6259, A2 => mult_143_n6078, ZN => 
                           mult_143_n6260);
   U131 : OAI21_X1 port map( B1 => n891, B2 => n882, A => n886, ZN => 
                           mult_143_n6078);
   U138 : AOI21_X1 port map( B1 => mult_143_n6605, B2 => n3803, A => n2707, ZN 
                           => mult_143_n5712);
   U142 : AND2_X1 port map( A1 => n3678, A2 => n971, ZN => n546);
   U144 : NAND2_X1 port map( A1 => n2906, A2 => B_SIG(16), ZN => n426);
   U145 : AOI22_X1 port map( A1 => B_SIG(7), A2 => n765, B1 => B_SIG(6), B2 => 
                           n787, ZN => mult_143_n6212);
   U147 : OAI22_X1 port map( A1 => n560, A2 => mult_143_n5705, B1 => n2869, B2 
                           => n4878, ZN => mult_143_n5709);
   U153 : XNOR2_X1 port map( A => mult_143_n5680, B => mult_143_n5679, ZN => 
                           n606);
   U157 : INV_X1 port map( A => B_SIG(23), ZN => n557);
   U165 : AND2_X1 port map( A1 => n3531, A2 => n4736, ZN => n508);
   U167 : OAI22_X1 port map( A1 => n812, A2 => n490, B1 => n825, B2 => n487, ZN
                           => mult_143_n6245);
   U174 : OAI21_X1 port map( B1 => mult_143_n6627, B2 => mult_143_n4842, A => 
                           mult_143_n5197, ZN => mult_143_n5196);
   U175 : AOI222_X1 port map( A1 => mult_143_n5598, A2 => mult_143_n5597, B1 =>
                           mult_143_n5598, B2 => n2846, C1 => mult_143_n5597, 
                           C2 => mult_143_n5596, ZN => mult_143_n5580);
   U179 : AND2_X1 port map( A1 => n3806, A2 => n4845, ZN => n395);
   U181 : XNOR2_X1 port map( A => A_SIG(21), B => A_SIG(22), ZN => 
                           mult_143_n6111);
   U186 : NOR2_X1 port map( A1 => B_SIG(18), A2 => B_SIG(17), ZN => 
                           mult_143_n6003);
   U188 : AND2_X1 port map( A1 => n3772, A2 => n3787, ZN => n436);
   U190 : AND2_X1 port map( A1 => n3798, A2 => n3788, ZN => n442);
   U196 : AOI21_X1 port map( B1 => mult_143_n48, B2 => B_SIG(7), A => 
                           mult_143_n6240, ZN => mult_143_n6239);
   U198 : OAI21_X1 port map( B1 => mult_143_n5580, B2 => n417, A => n416, ZN =>
                           n1508);
   U199 : AOI21_X1 port map( B1 => B_SIG(9), B2 => n1027, A => mult_143_n5196, 
                           ZN => mult_143_n5195);
   U202 : AOI21_X1 port map( B1 => B_SIG(7), B2 => mult_143_n6621, A => 
                           mult_143_n4819, ZN => mult_143_n4818);
   U203 : XNOR2_X1 port map( A => n1051, B => n4947, ZN => n1577);
   U204 : NOR2_X1 port map( A1 => mult_143_n4953, A2 => n395, ZN => n394);
   U207 : XNOR2_X1 port map( A => n1516, B => n4760, ZN => mult_143_n4991);
   U211 : NAND2_X1 port map( A1 => A_SIG(0), A2 => mult_143_n5853, ZN => 
                           mult_143_n5124);
   U215 : XNOR2_X1 port map( A => n532, B => n4750, ZN => n1574);
   U218 : AOI21_X1 port map( B1 => n4595, B2 => n4733, A => n1078, ZN => 
                           mult_143_n4903);
   U219 : AOI21_X1 port map( B1 => B_SIG(7), B2 => mult_143_n36, A => 
                           mult_143_n6193, ZN => mult_143_n6192);
   U229 : XNOR2_X1 port map( A => n3592, B => n1578, ZN => mult_143_n5232);
   U230 : AOI21_X1 port map( B1 => n4688, B2 => n3809, A => mult_143_n5903, ZN 
                           => n1507);
   U231 : XNOR2_X1 port map( A => n1559, B => n3739, ZN => mult_143_n5578);
   U233 : AOI222_X1 port map( A1 => n3496, A2 => n3702, B1 => n3739, B2 => 
                           n3496, C1 => n3739, C2 => n3702, ZN => n1473);
   U235 : XNOR2_X1 port map( A => mult_143_n5414, B => n3754, ZN => 
                           mult_143_n5209);
   U238 : OAI21_X1 port map( B1 => n3830, B2 => n548, A => n547, ZN => 
                           mult_143_n5187);
   U241 : AOI21_X1 port map( B1 => n3785, B2 => n3809, A => n3562, ZN => 
                           mult_143_n5899);
   U244 : OAI21_X1 port map( B1 => n3673, B2 => n1584, A => n3060, ZN => 
                           mult_143_n5959);
   U245 : AOI21_X1 port map( B1 => n3819, B2 => n3804, A => n1527, ZN => 
                           mult_143_n6043);
   U249 : OAI21_X1 port map( B1 => n3659, B2 => n1584, A => n3053, ZN => 
                           mult_143_n5854);
   U250 : NOR2_X1 port map( A1 => n948, A2 => mult_143_n5432, ZN => 
                           mult_143_n5430);
   U251 : XNOR2_X1 port map( A => n3773, B => n3553, ZN => n1573);
   U258 : XNOR2_X1 port map( A => n4754, B => mult_143_n4903, ZN => n1572);
   U259 : OAI21_X1 port map( B1 => n3792, B2 => n3791, A => mult_143_n4344, ZN 
                           => mult_143_n5191);
   U261 : XNOR2_X1 port map( A => n748, B => mult_143_n5230, ZN => n1571);
   U264 : XNOR2_X1 port map( A => mult_143_n5023, B => mult_143_n4490, ZN => 
                           mult_143_n5019);
   U274 : XNOR2_X1 port map( A => n445, B => n4657, ZN => mult_143_n1719);
   U277 : NAND2_X1 port map( A1 => mult_143_n5142, A2 => n1473, ZN => 
                           mult_143_n3083);
   U278 : NOR2_X1 port map( A1 => mult_143_n5142, A2 => n1473, ZN => n951);
   U300 : OAI21_X1 port map( B1 => mult_143_n6501, B2 => n951, A => 
                           mult_143_n3083, ZN => mult_143_n405);
   U302 : XNOR2_X1 port map( A => mult_143_n4928, B => n1626, ZN => n957);
   U304 : AOI21_X1 port map( B1 => mult_143_n3055, B2 => n1056, A => 
                           mult_143_n335, ZN => n1057);
   U306 : OR2_X1 port map( A1 => mult_143_n6124, A2 => n599, ZN => n1034);
   U307 : XNOR2_X1 port map( A => mult_143_n5999, B => B_SIG(19), ZN => n1035);
   U314 : INV_X1 port map( A => A_SIG(14), ZN => n649);
   U320 : INV_X1 port map( A => B_SIG(8), ZN => n886);
   U323 : OR2_X1 port map( A1 => mult_143_n5239, A2 => n4573, ZN => n1037);
   U324 : AND2_X1 port map( A1 => n1056, A2 => n1055, ZN => n1038);
   U329 : AND2_X1 port map( A1 => n391, A2 => n388, ZN => n1046);
   U332 : AOI21_X1 port map( B1 => B_SIG(15), B2 => B_SIG(17), A => B_SIG(16), 
                           ZN => mult_143_n6124);
   U333 : AND2_X1 port map( A1 => mult_143_n5300, A2 => n523, ZN => n1048);
   U337 : INV_X1 port map( A => B_SIG(9), ZN => n882);
   U341 : INV_X1 port map( A => B_SIG(7), ZN => n891);
   U346 : OR2_X1 port map( A1 => mult_143_n6198, A2 => n641, ZN => n1053);
   U350 : INV_X1 port map( A => mult_143_n4824, ZN => n382);
   U351 : INV_X1 port map( A => B_SIG(21), ZN => n847);
   U352 : OR2_X1 port map( A1 => mult_143_n6243, A2 => mult_143_n6244, ZN => 
                           n981);
   U354 : INV_X1 port map( A => B_SIG(16), ZN => n860);
   U355 : INV_X1 port map( A => B_SIG(6), ZN => n895);
   U365 : INV_X1 port map( A => B_SIG(10), ZN => n878);
   U370 : INV_X1 port map( A => B_SIG(19), ZN => n852);
   U374 : AOI222_X1 port map( A1 => n3745, A2 => n3660, B1 => n3745, B2 => 
                           n3497, C1 => n3660, C2 => n3497, ZN => 
                           mult_143_n5190);
   U390 : NOR2_X1 port map( A1 => mult_143_n2755, A2 => mult_143_n5434, ZN => 
                           n511);
   U393 : OAI21_X1 port map( B1 => n4663, B2 => mult_143_n373, A => 
                           mult_143_n5170, ZN => mult_143_n364);
   U394 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => mult_143_n4842, A => 
                           mult_143_n4888, ZN => mult_143_n4887);
   U395 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => mult_143_n4848, A => 
                           mult_143_n6194, ZN => mult_143_n6193);
   U396 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => mult_143_n4824, A => 
                           n486, ZN => n485);
   U398 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => mult_143_n4828, A => 
                           mult_143_n6241, ZN => mult_143_n6240);
   U402 : OR2_X1 port map( A1 => n2922, A2 => mult_143_n4768, ZN => n620);
   U403 : XNOR2_X1 port map( A => n2749, B => n3543, ZN => mult_143_n5004);
   U404 : NOR2_X1 port map( A1 => mult_143_n6115, A2 => n2825, ZN => n1060);
   U406 : NAND2_X1 port map( A1 => n4936, A2 => n2936, ZN => mult_143_n4789);
   U407 : XNOR2_X1 port map( A => mult_143_n5969, B => B_SIG(11), ZN => n1061);
   U410 : XNOR2_X1 port map( A => mult_143_n5969, B => B_SIG(11), ZN => 
                           mult_143_n3007);
   U412 : AOI21_X1 port map( B1 => n4714, B2 => n3820, A => mult_143_n6100, ZN 
                           => mult_143_n6099);
   U418 : AOI21_X1 port map( B1 => n3806, B2 => n4714, A => mult_143_n6064, ZN 
                           => mult_143_n6063);
   U419 : AOI21_X1 port map( B1 => n4626, B2 => n4672, A => n500, ZN => 
                           mult_143_n5052);
   U422 : AOI21_X1 port map( B1 => n3778, B2 => n3806, A => mult_143_n4923, ZN 
                           => mult_143_n4922);
   U423 : AOI21_X1 port map( B1 => n1062, B2 => n382, A => n456, ZN => n1505);
   U424 : XOR2_X1 port map( A => mult_143_n6102, B => mult_143_n6103, Z => 
                           n1062);
   U426 : AOI222_X1 port map( A1 => n1645, A2 => n3751, B1 => n1645, B2 => 
                           n3524, C1 => n3751, C2 => n3524, ZN => 
                           mult_143_n5441);
   U427 : AOI21_X1 port map( B1 => n2923, B2 => n2786, A => mult_143_n6578, ZN 
                           => n1063);
   U429 : AOI21_X1 port map( B1 => n774, B2 => B_SIG(10), A => mult_143_n4877, 
                           ZN => mult_143_n4876);
   U518 : XNOR2_X1 port map( A => mult_143_n5739, B => n3737, ZN => n1064);
   U557 : XNOR2_X1 port map( A => n3663, B => n3721, ZN => n1065);
   U564 : AOI222_X1 port map( A1 => n1049, A2 => mult_143_n5587, B1 => n1049, 
                           B2 => mult_143_n5588, C1 => mult_143_n5587, C2 => 
                           mult_143_n5588, ZN => n1067);
   U643 : XNOR2_X1 port map( A => B_SIG(5), B => mult_143_n6307, ZN => 
                           mult_143_n3096);
   U645 : XNOR2_X1 port map( A => B_SIG(5), B => mult_143_n6307, ZN => n1068);
   U648 : OAI22_X1 port map( A1 => mult_143_n5667, A2 => n546, B1 => n3678, B2 
                           => n971, ZN => mult_143_n5658);
   U649 : NAND2_X1 port map( A1 => mult_143_n6079, A2 => mult_143_n6260, ZN => 
                           n1069);
   U651 : XNOR2_X1 port map( A => mult_143_n5638, B => n3631, ZN => 
                           mult_143_n5625);
   U652 : AOI222_X1 port map( A1 => n4874, A2 => mult_143_n5616, B1 => 
                           mult_143_n5615, B2 => n4875, C1 => mult_143_n5617, 
                           C2 => mult_143_n5616, ZN => mult_143_n5426);
   U655 : OAI21_X1 port map( B1 => mult_143_n5439, B2 => n1064, A => n953, ZN 
                           => mult_143_n3448);
   U656 : AOI21_X1 port map( B1 => n2908, B2 => n3817, A => mult_143_n4901, ZN 
                           => mult_143_n4900);
   U657 : OAI22_X1 port map( A1 => mult_143_n4896, A2 => n482, B1 => n4630, B2 
                           => n1572, ZN => mult_143_n897);
   U658 : XNOR2_X1 port map( A => mult_143_n4900, B => n4625, ZN => 
                           mult_143_n4896);
   U659 : AND2_X1 port map( A1 => n480, A2 => n479, ZN => mult_143_n6113);
   U667 : AOI222_X1 port map( A1 => n3690, A2 => n3559, B1 => n3690, B2 => 
                           n1573, C1 => n3559, C2 => n1573, ZN => mult_143_n977
                           );
   U670 : AOI21_X1 port map( B1 => B_SIG(10), B2 => n799, A => mult_143_n4960, 
                           ZN => mult_143_n4959);
   U672 : NAND2_X1 port map( A1 => mult_143_n5467, A2 => n515, ZN => n514);
   U674 : NOR2_X1 port map( A1 => mult_143_n5446, A2 => mult_143_n5445, ZN => 
                           mult_143_n2755);
   U676 : INV_X1 port map( A => mult_143_n5758, ZN => n698);
   U686 : XNOR2_X1 port map( A => n1575, B => n3493, ZN => mult_143_n5754);
   U698 : XNOR2_X1 port map( A => n493, B => n2840, ZN => n1568);
   U701 : NOR2_X1 port map( A1 => mult_143_n5033, A2 => n494, ZN => n493);
   U702 : AOI21_X1 port map( B1 => n2908, B2 => n4665, A => mult_143_n6005, ZN 
                           => mult_143_n6004);
   U720 : AOI21_X1 port map( B1 => n2908, B2 => n3809, A => mult_143_n5906, ZN 
                           => mult_143_n5905);
   U721 : AND2_X1 port map( A1 => n1563, A2 => n4625, ZN => n558);
   U724 : OAI22_X1 port map( A1 => n558, A2 => mult_143_n4972, B1 => n4625, B2 
                           => n1563, ZN => mult_143_n809);
   U726 : OAI21_X1 port map( B1 => mult_143_n6625, B2 => mult_143_n4820, A => 
                           mult_143_n5194, ZN => mult_143_n5193);
   U729 : XNOR2_X1 port map( A => mult_143_n6035, B => B_SIG(15), ZN => 
                           mult_143_n6625);
   U730 : XNOR2_X1 port map( A => n568, B => n1839, ZN => n1567);
   U731 : XNOR2_X1 port map( A => mult_143_n6112, B => n557, ZN => n1071);
   U732 : XNOR2_X1 port map( A => mult_143_n5089, B => n4752, ZN => n660);
   U735 : XNOR2_X1 port map( A => n441, B => n4754, ZN => mult_143_n4972);
   U736 : INV_X1 port map( A => n1072, ZN => mult_143_n6031);
   U744 : AOI21_X1 port map( B1 => n4871, B2 => n3801, A => mult_143_n5845, ZN 
                           => mult_143_n5844);
   U754 : XNOR2_X1 port map( A => n1600, B => n2780, ZN => mult_143_n5035);
   U756 : INV_X1 port map( A => n433, ZN => n532);
   U757 : XNOR2_X1 port map( A => n424, B => n423, ZN => n1565);
   U762 : XNOR2_X1 port map( A => n424, B => n423, ZN => n1075);
   U767 : XNOR2_X1 port map( A => n424, B => n423, ZN => mult_143_n6624);
   U769 : OAI21_X1 port map( B1 => mult_143_n5970, B2 => n539, A => n537, ZN =>
                           mult_143_n5969);
   U773 : AOI21_X1 port map( B1 => n3804, B2 => n3817, A => n1526, ZN => 
                           mult_143_n5956);
   U774 : INV_X1 port map( A => mult_143_n5426, ZN => n724);
   U775 : AOI222_X1 port map( A1 => n3504, A2 => n4590, B1 => n3504, B2 => 
                           mult_143_n4965, C1 => n4590, C2 => mult_143_n4965, 
                           ZN => mult_143_n811);
   U776 : XNOR2_X1 port map( A => n649, B => mult_143_n4818, ZN => n1564);
   U777 : XNOR2_X1 port map( A => n527, B => n3773, ZN => n1563);
   U780 : NOR2_X1 port map( A1 => mult_143_n4980, A2 => n528, ZN => n527);
   U781 : OAI21_X1 port map( B1 => mult_143_n4757, B2 => mult_143_n6498, A => 
                           n944, ZN => mult_143_n4755);
   U784 : AOI21_X1 port map( B1 => mult_143_n4755, B2 => n2764, A => 
                           mult_143_n6499, ZN => n385);
   U785 : AOI222_X1 port map( A1 => mult_143_n4984, A2 => n4670, B1 => 
                           mult_143_n4984, B2 => n4579, C1 => mult_143_n6367, 
                           C2 => n4579, ZN => mult_143_n795);
   U808 : AOI222_X1 port map( A1 => n4720, A2 => mult_143_n5186, B1 => n4720, 
                           B2 => n2909, C1 => n2909, C2 => mult_143_n5186, ZN 
                           => n1470);
   U812 : INV_X1 port map( A => mult_143_n5695, ZN => n745);
   U813 : AOI22_X1 port map( A1 => mult_143_n6597, A2 => n745, B1 => 
                           mult_143_n5695, B2 => n4650, ZN => mult_143_n5694);
   U815 : NAND2_X1 port map( A1 => mult_143_n5189, A2 => mult_143_n5190, ZN => 
                           mult_143_n4502);
   U817 : XNOR2_X1 port map( A => n1501, B => n4754, ZN => mult_143_n4869);
   U819 : AOI21_X1 port map( B1 => n3786, B2 => n3802, A => n3561, ZN => n1503)
                           ;
   U824 : AOI21_X1 port map( B1 => n4890, B2 => n3802, A => mult_143_n4874, ZN 
                           => n1501);
   U825 : AOI21_X1 port map( B1 => n2908, B2 => n3802, A => mult_143_n4920, ZN 
                           => mult_143_n4919);
   U826 : NAND2_X1 port map( A1 => n3802, A2 => n4695, ZN => n1079);
   U827 : AOI22_X1 port map( A1 => B_SIG(9), A2 => n765, B1 => B_SIG(8), B2 => 
                           n787, ZN => mult_143_n6241);
   U829 : AOI222_X1 port map( A1 => n1567, A2 => mult_143_n4994, B1 => 
                           mult_143_n4994, B2 => n4580, C1 => n1567, C2 => 
                           n4580, ZN => mult_143_n777);
   U835 : OAI21_X1 port map( B1 => mult_143_n4891, B2 => mult_143_n3010, A => 
                           mult_143_n5002, ZN => mult_143_n5001);
   U842 : OAI221_X1 port map( B1 => mult_143_n6125, B2 => n1069, C1 => 
                           mult_143_n6125, C2 => mult_143_n6127, A => 
                           mult_143_n6128, ZN => n1077);
   U860 : NAND2_X1 port map( A1 => mult_143_n5440, A2 => mult_143_n5441, ZN => 
                           n953);
   U861 : OAI21_X1 port map( B1 => mult_143_n6628, B2 => mult_143_n4820, A => 
                           mult_143_n4821, ZN => mult_143_n4819);
   U862 : AOI21_X1 port map( B1 => n4890, B2 => n3823, A => mult_143_n4857, ZN 
                           => mult_143_n4856);
   U869 : XNOR2_X1 port map( A => mult_143_n5069, B => n1839, ZN => 
                           mult_143_n5067);
   U870 : XNOR2_X1 port map( A => n3648, B => n1839, ZN => n1560);
   U875 : AOI21_X1 port map( B1 => n1035, B2 => n382, A => n380, ZN => n1500);
   U877 : XNOR2_X1 port map( A => mult_143_n5004, B => n3792, ZN => n972);
   U878 : OAI21_X1 port map( B1 => mult_143_n3137, B2 => mult_143_n4820, A => 
                           mult_143_n4943, ZN => mult_143_n4942);
   U880 : OAI21_X1 port map( B1 => n3666, B2 => n3596, A => mult_143_n5444, ZN 
                           => mult_143_n5443);
   U884 : XNOR2_X1 port map( A => mult_143_n4937, B => n3791, ZN => n608);
   U886 : XNOR2_X1 port map( A => mult_143_n4941, B => n3773, ZN => 
                           mult_143_n4937);
   U890 : OAI22_X1 port map( A1 => mult_143_n6630, A2 => mult_143_n4891, B1 => 
                           n910, B2 => n982, ZN => mult_143_n5231);
   U893 : OAI21_X1 port map( B1 => mult_143_n6630, B2 => mult_143_n4842, A => 
                           mult_143_n4843, ZN => mult_143_n4841);
   U894 : INV_X1 port map( A => mult_143_n5228, ZN => n671);
   U897 : NOR2_X1 port map( A1 => mult_143_n5939, A2 => mult_143_n6029, ZN => 
                           mult_143_n6028);
   U899 : AOI222_X1 port map( A1 => mult_143_n5760, A2 => n4673, B1 => n4653, 
                           B2 => mult_143_n5760, C1 => n3101, C2 => n4673, ZN 
                           => n1469);
   U900 : XNOR2_X1 port map( A => mult_143_n5456, B => n3650, ZN => 
                           mult_143_n5445);
   U901 : XNOR2_X1 port map( A => n4653, B => mult_143_n5769, ZN => n1558);
   U902 : NAND2_X1 port map( A1 => mult_143_n4905, A2 => n1079, ZN => n1078);
   U906 : XNOR2_X1 port map( A => n1083, B => n2686, ZN => n992);
   U907 : XNOR2_X1 port map( A => n3690, B => n3559, ZN => n1083);
   U908 : XNOR2_X1 port map( A => mult_143_n5999, B => n852, ZN => n1085);
   U911 : OAI21_X1 port map( B1 => n3596, B2 => n3667, A => mult_143_n4927, ZN 
                           => mult_143_n4926);
   U913 : OAI21_X1 port map( B1 => n3594, B2 => n3667, A => mult_143_n4881, ZN 
                           => mult_143_n4880);
   U915 : OAI21_X1 port map( B1 => n3667, B2 => n3644, A => mult_143_n4864, ZN 
                           => mult_143_n4863);
   U918 : NOR2_X1 port map( A1 => mult_143_n5027, A2 => n572, ZN => n571);
   U919 : AOI21_X1 port map( B1 => n637, B2 => B_SIG(15), A => mult_143_n6085, 
                           ZN => n425);
   U920 : OAI21_X1 port map( B1 => n637, B2 => n1034, A => mult_143_n6106, ZN 
                           => n480);
   U922 : XNOR2_X1 port map( A => n3627, B => n3815, ZN => mult_143_n5638);
   U925 : AOI22_X1 port map( A1 => mult_143_n1530, A2 => n1556, B1 => n2690, B2
                           => mult_143_n1901, ZN => mult_143_n724);
   U933 : XNOR2_X1 port map( A => n507, B => n2840, ZN => n1556);
   U934 : NOR2_X1 port map( A1 => mult_143_n5046, A2 => n508, ZN => n507);
   U935 : OR2_X1 port map( A1 => mult_143_n5187, A2 => mult_143_n5188, ZN => 
                           n604);
   U936 : AND2_X1 port map( A1 => mult_143_n5188, A2 => mult_143_n5187, ZN => 
                           n605);
   U939 : AOI21_X1 port map( B1 => n772, B2 => B_SIG(17), A => mult_143_n4970, 
                           ZN => n1499);
   U953 : XNOR2_X1 port map( A => n607, B => B_SIG(21), ZN => n1555);
   U979 : OAI21_X1 port map( B1 => n563, B2 => mult_143_n5724, A => n562, ZN =>
                           mult_143_n5733);
   U982 : AOI222_X1 port map( A1 => mult_143_n5709, A2 => mult_143_n5707, B1 =>
                           mult_143_n5709, B2 => mult_143_n5708, C1 => 
                           mult_143_n5707, C2 => mult_143_n5708, ZN => 
                           mult_143_n5724);
   U984 : OR2_X1 port map( A1 => mult_143_n5206, A2 => mult_143_n5207, ZN => 
                           n942);
   U985 : INV_X1 port map( A => n1055, ZN => mult_143_n4340);
   U990 : INV_X1 port map( A => n1039, ZN => mult_143_n6513);
   U995 : INV_X1 port map( A => mult_143_n522, ZN => n1718);
   U1003 : INV_X1 port map( A => n1056, ZN => mult_143_n6518);
   U1010 : INV_X1 port map( A => mult_143_n904, ZN => n1722);
   U1015 : INV_X1 port map( A => mult_143_n744, ZN => mult_143_n6361);
   U1037 : INV_X1 port map( A => mult_143_n581, ZN => mult_143_n6309);
   U1038 : INV_X1 port map( A => mult_143_n922, ZN => n1723);
   U1045 : INV_X1 port map( A => mult_143_n938, ZN => n1728);
   U1046 : INV_X1 port map( A => mult_143_n3455, ZN => mult_143_n6570);
   U1063 : INV_X1 port map( A => n1040, ZN => mult_143_n6379);
   U1102 : INV_X1 port map( A => n1042, ZN => mult_143_n6573);
   U1111 : INV_X1 port map( A => n945, ZN => mult_143_n6499);
   U1112 : INV_X1 port map( A => n4731, ZN => mult_143_n6510);
   U1113 : INV_X1 port map( A => n954, ZN => mult_143_n6559);
   U1114 : INV_X1 port map( A => n944, ZN => mult_143_n4351);
   U1116 : INV_X1 port map( A => n953, ZN => mult_143_n6523);
   U1118 : INV_X1 port map( A => n948, ZN => mult_143_n4357);
   U1119 : INV_X1 port map( A => n949, ZN => mult_143_n4363);
   U1120 : INV_X1 port map( A => n951, ZN => mult_143_n4348);
   U1121 : INV_X1 port map( A => n971, ZN => mult_143_n6598);
   U1122 : INV_X1 port map( A => n967, ZN => mult_143_n6406);
   U1147 : INV_X1 port map( A => mult_143_n795, ZN => mult_143_n6368);
   U1154 : INV_X1 port map( A => n1047, ZN => mult_143_n6532);
   U1163 : INV_X1 port map( A => n4870, ZN => mult_143_n4475);
   U1164 : INV_X1 port map( A => n1045, ZN => mult_143_n6397);
   U1181 : INV_X1 port map( A => n4892, ZN => mult_143_n6580);
   U1199 : INV_X1 port map( A => n4728, ZN => mult_143_n4359);
   U1201 : INV_X1 port map( A => mult_143_n6620, ZN => mult_143_n6491);
   U1205 : INV_X1 port map( A => mult_143_n3075, ZN => mult_143_n6535);
   U1207 : INV_X1 port map( A => mult_143_n344, ZN => mult_143_n4339);
   U1210 : INV_X1 port map( A => mult_143_n304, ZN => mult_143_n4366);
   U1212 : INV_X1 port map( A => mult_143_n4502, ZN => mult_143_n6526);
   U1213 : INV_X1 port map( A => n2891, ZN => mult_143_n6490);
   U1225 : INV_X1 port map( A => mult_143_n4344, ZN => mult_143_n6473);
   U1228 : INV_X1 port map( A => mult_143_n1719, ZN => mult_143_n6610);
   U1232 : INV_X1 port map( A => mult_143_n1753, ZN => mult_143_n4361);
   U1233 : INV_X1 port map( A => mult_143_n4493, ZN => mult_143_n6516);
   U1235 : INV_X1 port map( A => mult_143_n412, ZN => mult_143_n6501);
   U1237 : INV_X1 port map( A => mult_143_n1059, ZN => mult_143_n6478);
   U1242 : INV_X1 port map( A => n419, ZN => mult_143_n6607);
   U1244 : INV_X1 port map( A => n4887, ZN => mult_143_n6517);
   U1245 : INV_X1 port map( A => mult_143_n373, ZN => mult_143_n6536);
   U1253 : INV_X1 port map( A => mult_143_n218, ZN => mult_143_n6524);
   U1277 : INV_X1 port map( A => A_EXP(7), ZN => n25);
   U1278 : INV_X1 port map( A => B_EXP(7), ZN => n24);
   U1284 : INV_X1 port map( A => n992, ZN => mult_143_n6407);
   U1285 : INV_X1 port map( A => n957, ZN => mult_143_n6374);
   U1291 : INV_X1 port map( A => n991, ZN => mult_143_n4355);
   U1293 : INV_X1 port map( A => n965, ZN => mult_143_n6564);
   U1294 : INV_X1 port map( A => n968, ZN => mult_143_n6388);
   U1307 : INV_X1 port map( A => mult_143_n276, ZN => mult_143_n6578);
   U1311 : INV_X1 port map( A => n972, ZN => mult_143_n6551);
   U1312 : INV_X1 port map( A => n963, ZN => mult_143_n6549);
   U1316 : INV_X1 port map( A => mult_143_n1116, ZN => n1759);
   U1317 : INV_X1 port map( A => mult_143_n364, ZN => mult_143_n6550);
   U1223 : INV_X1 port map( A => mult_143_n813, ZN => mult_143_n6592);
   U1276 : INV_X1 port map( A => mult_143_n1754, ZN => mult_143_n6408);
   U1215 : INV_X1 port map( A => mult_143_n759, ZN => mult_143_n6362);
   U1136 : INV_X1 port map( A => mult_143_n809, ZN => mult_143_n6589);
   U1287 : INV_X1 port map( A => n970, ZN => mult_143_n6543);
   U1318 : INV_X1 port map( A => n969, ZN => mult_143_n6369);
   mult_143_U4660 : XOR2_X1 port map( A => A_SIG(7), B => A_SIG(8), Z => 
                           mult_143_n6253);
   mult_143_U4671 : XOR2_X1 port map( A => A_SIG(20), B => A_SIG(19), Z => 
                           mult_143_n6300);
   U558 : INV_X1 port map( A => mult_143_n6244, ZN => n646);
   U727 : NOR2_X1 port map( A1 => mult_143_n6300, A2 => mult_143_n6293, ZN => 
                           mult_143_n74);
   U795 : AND3_X1 port map( A1 => mult_143_n6300, A2 => mult_143_n6293, A3 => 
                           mult_143_n6301, ZN => mult_143_n84);
   U51 : AND3_X1 port map( A1 => mult_143_n6284, A2 => mult_143_n6181, A3 => 
                           mult_143_n6292, ZN => mult_143_n6621);
   U208 : CLKBUF_X1 port map( A => mult_143_n74, Z => n778);
   U140 : OAI211_X1 port map( C1 => B_SIG(14), C2 => B_SIG(15), A => 
                           mult_143_n6030, B => n636, ZN => mult_143_n6125);
   U90 : INV_X1 port map( A => n980, ZN => n1031);
   mult_143_U3934 : AND3_X1 port map( A1 => mult_143_n6243, A2 => 
                           mult_143_n6244, A3 => mult_143_n6242, ZN => 
                           mult_143_n48);
   U821 : NAND2_X1 port map( A1 => n646, A2 => mult_143_n6243, ZN => 
                           mult_143_n4828);
   U1177 : INV_X1 port map( A => mult_143_n901, ZN => mult_143_n6382);
   U1175 : INV_X1 port map( A => mult_143_n886, ZN => mult_143_n6541);
   U81 : INV_X1 port map( A => n1053, ZN => n1026);
   U431 : INV_X1 port map( A => n1052, ZN => n787);
   U1131 : INV_X1 port map( A => mult_143_n724, ZN => mult_143_n6360);
   U1206 : INV_X1 port map( A => mult_143_n3073, ZN => mult_143_n6498);
   U1191 : INV_X1 port map( A => n1050, ZN => mult_143_n6398);
   U32 : AOI222_X1 port map( A1 => n2837, A2 => n4863, B1 => n2837, B2 => 
                           mult_143_n6401, C1 => n4863, C2 => mult_143_n6401, 
                           ZN => mult_143_n5598);
   U50 : INV_X1 port map( A => n996, ZN => n2599);
   U53 : AOI222_X1 port map( A1 => n4585, A2 => n2750, B1 => n4585, B2 => n3831
                           , C1 => n2750, C2 => n3831, ZN => mult_143_n5660);
   U80 : NOR2_X1 port map( A1 => n3005, A2 => mult_143_n335, ZN => n3004);
   U103 : XNOR2_X1 port map( A => n3029, B => mult_143_n5020, ZN => n2869);
   U104 : AOI21_X1 port map( B1 => n3029, B2 => n2716, A => n3028, ZN => 
                           mult_143_n6554);
   U106 : OAI22_X1 port map( A1 => mult_143_n4948, A2 => n2720, B1 => n4590, B2
                           => n4630, ZN => n969);
   U107 : AOI21_X1 port map( B1 => n2803, B2 => mult_143_n6432, A => 
                           mult_143_n6434, ZN => n2994);
   U124 : XNOR2_X1 port map( A => n2755, B => n2959, ZN => mult_143_n5725);
   U125 : OAI22_X1 port map( A1 => mult_143_n4852, A2 => n3001, B1 => n1590, B2
                           => n1614, ZN => n1050);
   U128 : NOR2_X1 port map( A1 => mult_143_n6061, A2 => n2986, ZN => n2985);
   U135 : XNOR2_X1 port map( A => mult_143_n5887, B => n3099, ZN => 
                           mult_143_n6434);
   U137 : AND2_X1 port map( A1 => mult_143_n6272, A2 => n2976, ZN => n632);
   U139 : XNOR2_X1 port map( A => n2804, B => n3686, ZN => n2803);
   U141 : NOR2_X1 port map( A1 => n3040, A2 => n3039, ZN => mult_143_n706);
   U151 : NAND2_X1 port map( A1 => n654, A2 => mult_143_n6110, ZN => 
                           mult_143_n4891);
   U152 : XNOR2_X1 port map( A => n2988, B => n4570, ZN => mult_143_n5153);
   U158 : OR2_X1 port map( A1 => n2793, A2 => n2792, ZN => n2791);
   U172 : INV_X1 port map( A => mult_143_n2772, ZN => n2600);
   U178 : NOR2_X1 port map( A1 => n4768, A2 => n1560, ZN => n3028);
   U191 : OAI21_X1 port map( B1 => n4619, B2 => n4621, A => n4584, ZN => n2865)
                           ;
   U213 : AND2_X1 port map( A1 => n3494, A2 => n3705, ZN => mult_143_n5641);
   U214 : AND2_X1 port map( A1 => n3806, A2 => n3784, ZN => n2986);
   U224 : NAND2_X1 port map( A1 => n2841, A2 => n2971, ZN => mult_143_n6030);
   U254 : INV_X1 port map( A => A_SIG(8), ZN => n1782);
   U256 : XNOR2_X1 port map( A => A_SIG(8), B => A_SIG(9), ZN => mult_143_n6244
                           );
   U257 : AND2_X1 port map( A1 => n3817, A2 => n3780, ZN => n2958);
   U265 : NOR2_X1 port map( A1 => n3756, A2 => n3548, ZN => n2792);
   U266 : NOR2_X1 port map( A1 => mult_143_n6518, A2 => mult_143_n4475, ZN => 
                           n3005);
   U267 : NOR2_X1 port map( A1 => n2978, A2 => B_SIG(6), ZN => n2974);
   U269 : AOI21_X1 port map( B1 => mult_143_n5058, B2 => n3824, A => 
                           mult_143_n1900, ZN => n3040);
   U273 : OR2_X1 port map( A1 => n442, A2 => n2952, ZN => n2951);
   U279 : AND2_X1 port map( A1 => n3510, A2 => n3742, ZN => n2794);
   U282 : INV_X1 port map( A => mult_143_n5439, ZN => n2920);
   U283 : INV_X1 port map( A => mult_143_n1039, ZN => mult_143_n6432);
   U291 : INV_X1 port map( A => mult_143_n1005, ZN => mult_143_n6417);
   U299 : AOI222_X1 port map( A1 => B_SIG(14), A2 => B_SIG(15), B1 => B_SIG(14)
                           , B2 => mult_143_n6129, C1 => mult_143_n6129, C2 => 
                           B_SIG(15), ZN => mult_143_n6128);
   U301 : NAND2_X1 port map( A1 => n632, A2 => n2974, ZN => n2973);
   U303 : XNOR2_X1 port map( A => n394, B => n1839, ZN => mult_143_n4948);
   U309 : NAND2_X1 port map( A1 => n2978, A2 => n2977, ZN => n2976);
   U311 : XNOR2_X1 port map( A => mult_143_n5145, B => n2782, ZN => 
                           mult_143_n5144);
   U322 : INV_X1 port map( A => n946, ZN => mult_143_n6560);
   U330 : XNOR2_X1 port map( A => mult_143_n4856, B => n4625, ZN => 
                           mult_143_n4852);
   U335 : INV_X1 port map( A => mult_143_n1027, ZN => mult_143_n6427);
   U348 : NOR2_X1 port map( A1 => B_SIG(13), A2 => B_SIG(14), ZN => 
                           mult_143_n6029);
   U353 : INV_X1 port map( A => mult_143_n671, ZN => mult_143_n6348);
   U357 : XNOR2_X1 port map( A => n2985, B => n4750, ZN => mult_143_n1582);
   U359 : INV_X1 port map( A => mult_143_n977, ZN => mult_143_n6402);
   U377 : NAND2_X1 port map( A1 => B_SIG(13), A2 => B_SIG(14), ZN => 
                           mult_143_n5940);
   U381 : XNOR2_X1 port map( A => n2606, B => n4632, ZN => n2959);
   U382 : INV_X1 port map( A => mult_143_n917, ZN => mult_143_n6385);
   U384 : XNOR2_X1 port map( A => mult_143_n706, B => n3042, ZN => 
                           mult_143_n5742);
   U397 : INV_X1 port map( A => mult_143_n610, ZN => mult_143_n6322);
   U415 : NOR2_X1 port map( A1 => mult_143_n1894, A2 => n2620, ZN => 
                           mult_143_n5543);
   U417 : XNOR2_X1 port map( A => A_SIG(20), B => A_SIG(21), ZN => 
                           mult_143_n4832);
   U449 : AOI21_X1 port map( B1 => n616, B2 => n1066, A => n2757, ZN => n1049);
   U472 : INV_X1 port map( A => mult_143_n897, ZN => mult_143_n6381);
   U504 : OR2_X1 port map( A1 => n646, A2 => mult_143_n6242, ZN => n1052);
   U511 : AND3_X1 port map( A1 => mult_143_n6253, A2 => mult_143_n6255, A3 => 
                           n643, ZN => mult_143_n36);
   U512 : AND3_X1 port map( A1 => mult_143_n6198, A2 => n641, A3 => 
                           mult_143_n6200, ZN => mult_143_n3228);
   U515 : INV_X1 port map( A => n981, ZN => n765);
   U529 : XOR2_X1 port map( A => mult_143_n5232, B => n3503, Z => n2601);
   U531 : AND2_X1 port map( A1 => mult_143_n412, A2 => n4724, ZN => n2602);
   U535 : AND2_X1 port map( A1 => mult_143_n3083, A2 => n4724, ZN => n2603);
   U543 : NOR2_X1 port map( A1 => mult_143_n5607, A2 => n2791, ZN => 
                           mult_143_n4493);
   U549 : AND2_X1 port map( A1 => mult_143_n5152, A2 => mult_143_n5153, ZN => 
                           n2604);
   U555 : OR2_X1 port map( A1 => n2690, A2 => mult_143_n1901, ZN => n2606);
   U560 : XNOR2_X1 port map( A => mult_143_n5847, B => n4670, ZN => n2608);
   U561 : XNOR2_X1 port map( A => n4670, B => mult_143_n5850, ZN => n2609);
   U584 : XOR2_X1 port map( A => n1064, B => mult_143_n5439, Z => n2611);
   U592 : INV_X1 port map( A => B_SIG(5), ZN => n2978);
   U596 : XOR2_X1 port map( A => n3674, B => n553, Z => n2612);
   U598 : XOR2_X1 port map( A => n3742, B => n3510, Z => n2614);
   U599 : XNOR2_X1 port map( A => n1632, B => n1588, ZN => n2615);
   U600 : INV_X1 port map( A => mult_143_n867, ZN => mult_143_n5666);
   U619 : NOR2_X1 port map( A1 => n2718, A2 => n4605, ZN => mult_143_n867);
   U624 : OR2_X1 port map( A1 => n2780, A2 => n2751, ZN => n2617);
   U626 : XNOR2_X1 port map( A => n4670, B => n1539, ZN => n2618);
   U627 : XNOR2_X1 port map( A => n1538, B => n3773, ZN => n2619);
   U628 : OR2_X1 port map( A1 => mult_143_n1895, A2 => n2731, ZN => n2620);
   U629 : XNOR2_X1 port map( A => mult_143_n6367, B => n1537, ZN => n2621);
   U630 : XNOR2_X1 port map( A => n3803, B => n1536, ZN => n2622);
   U632 : OR2_X1 port map( A1 => n4625, A2 => mult_143_n5035, ZN => n2624);
   U633 : OR2_X1 port map( A1 => mult_143_n5075, A2 => n4768, ZN => n2627);
   U644 : AND2_X1 port map( A1 => n2780, A2 => n4634, ZN => n2630);
   U647 : XOR2_X1 port map( A => n3741, B => n1665, Z => n2632);
   U653 : XNOR2_X1 port map( A => n2840, B => n1531, ZN => n2633);
   U654 : XNOR2_X1 port map( A => mult_143_n4490, B => n1530, ZN => n2634);
   U665 : OR2_X1 port map( A1 => mult_143_n6347, A2 => mult_143_n6348, ZN => 
                           n2636);
   U666 : AND2_X1 port map( A1 => mult_143_n5170, A2 => n4936, ZN => n2637);
   U687 : AND2_X1 port map( A1 => n744, A2 => mult_143_n5205, ZN => n2638);
   U719 : XOR2_X1 port map( A => mult_143_n6112, B => n557, Z => n1840);
   U733 : XNOR2_X1 port map( A => n536, B => mult_143_n5799, ZN => n1756);
   U737 : XNOR2_X1 port map( A => n536, B => mult_143_n5802, ZN => n1755);
   U739 : XNOR2_X1 port map( A => n536, B => mult_143_n5805, ZN => n1754);
   U740 : XNOR2_X1 port map( A => n3769, B => n3587, ZN => n1758);
   U748 : XNOR2_X1 port map( A => n3769, B => n3585, ZN => n1757);
   U750 : XNOR2_X1 port map( A => n642, B => mult_143_n5866, ZN => n1739);
   U751 : XNOR2_X1 port map( A => n642, B => mult_143_n5869, ZN => n1741);
   U763 : XNOR2_X1 port map( A => n642, B => mult_143_n5872, ZN => n1738);
   U764 : XNOR2_X1 port map( A => n642, B => mult_143_n5878, ZN => n1742);
   U765 : XNOR2_X1 port map( A => n3768, B => n3586, ZN => n1752);
   U766 : XNOR2_X1 port map( A => n1782, B => mult_143_n5920, ZN => n1719);
   U771 : XNOR2_X1 port map( A => n1782, B => mult_143_n5923, ZN => n1745);
   U779 : XOR2_X1 port map( A => A_SIG(20), B => mult_143_n6048, Z => n1730);
   U782 : XOR2_X1 port map( A => A_SIG(20), B => mult_143_n6054, Z => n1736);
   U786 : XOR2_X1 port map( A => A_SIG(20), B => mult_143_n6057, Z => n1734);
   U788 : XOR2_X1 port map( A => A_SIG(20), B => mult_143_n6051, Z => n1733);
   U791 : XOR2_X1 port map( A => mult_143_n4830, B => mult_143_n4831, Z => 
                           n1727);
   U793 : XOR2_X1 port map( A => n748, B => mult_143_n6068, Z => n1737);
   U794 : XOR2_X1 port map( A => n748, B => mult_143_n6071, Z => n1735);
   U798 : XOR2_X1 port map( A => mult_143_n5095, B => n2780, Z => n2664);
   U800 : OR2_X1 port map( A1 => n4670, A2 => mult_143_n1902, ZN => n2665);
   U809 : XNOR2_X1 port map( A => n1545, B => n3774, ZN => n2668);
   U810 : XNOR2_X1 port map( A => mult_143_n4490, B => n1543, ZN => n2669);
   U811 : XOR2_X1 port map( A => n4763, B => mult_143_n5187, Z => n2670);
   U820 : XNOR2_X1 port map( A => mult_143_n5814, B => n4670, ZN => n1749);
   U823 : XOR2_X1 port map( A => n1629, B => mult_143_n5015, Z => n2675);
   U830 : XNOR2_X1 port map( A => n4754, B => mult_143_n5966, ZN => n2679);
   U841 : XNOR2_X1 port map( A => n3822, B => n4768, ZN => n2692);
   U844 : OR2_X1 port map( A1 => n2685, A2 => n3803, ZN => n2694);
   U846 : XOR2_X1 port map( A => n4750, B => mult_143_n6063, Z => n2696);
   U847 : XOR2_X1 port map( A => A_SIG(17), B => mult_143_n6009, Z => n1729);
   U849 : OR2_X1 port map( A1 => n3803, A2 => n4586, ZN => n2704);
   U850 : XNOR2_X1 port map( A => mult_143_n6367, B => n1514, ZN => n2705);
   U854 : XNOR2_X1 port map( A => mult_143_n4490, B => mult_143_n6004, ZN => 
                           n2707);
   U855 : AND2_X1 port map( A1 => mult_143_n1815, A2 => n1765, ZN => n2709);
   U863 : AND2_X1 port map( A1 => mult_143_n6516, A2 => n4887, ZN => n2710);
   U864 : XNOR2_X1 port map( A => n4634, B => n2780, ZN => n2714);
   U866 : XOR2_X1 port map( A => mult_143_n5075, B => n3794, Z => n2715);
   U868 : NAND2_X1 port map( A1 => n1560, A2 => n4768, ZN => n2716);
   U872 : XOR2_X1 port map( A => mult_143_n5035, B => n3793, Z => n2717);
   U874 : OR2_X1 port map( A1 => mult_143_n5004, A2 => n4590, ZN => n2719);
   U879 : AND2_X1 port map( A1 => n4630, A2 => n4590, ZN => n2720);
   U882 : AND2_X1 port map( A1 => n3007, A2 => n3006, ZN => n2721);
   U888 : AND2_X1 port map( A1 => n3533, A2 => n3789, ZN => n2722);
   U896 : XOR2_X1 port map( A => n1664, B => mult_143_n6186, Z => n2723);
   U898 : XOR2_X1 port map( A => n3713, B => mult_143_n6162, Z => n2725);
   U909 : XNOR2_X1 port map( A => n2780, B => n2751, ZN => n2726);
   U910 : XNOR2_X1 port map( A => mult_143_n5956, B => n3803, ZN => n2727);
   U912 : XOR2_X1 port map( A => n1521, B => n473, Z => n2728);
   U917 : XOR2_X1 port map( A => n2840, B => mult_143_n6099, Z => n2731);
   U923 : XNOR2_X1 port map( A => n2840, B => mult_143_n6119, ZN => n2733);
   U927 : XNOR2_X1 port map( A => n3662, B => n3616, ZN => n2736);
   U928 : XOR2_X1 port map( A => n1623, B => mult_143_n4883, Z => n2737);
   U929 : XNOR2_X1 port map( A => n1529, B => n3792, ZN => n2739);
   U938 : XNOR2_X1 port map( A => mult_143_n6135, B => mult_143_n6136, ZN => 
                           n1725);
   U940 : XOR2_X1 port map( A => A_SIG(8), B => mult_143_n5918, Z => n1748);
   U941 : XOR2_X1 port map( A => A_SIG(8), B => mult_143_n5916, Z => n1740);
   U942 : XNOR2_X1 port map( A => mult_143_n6137, B => mult_143_n6138, ZN => 
                           n1720);
   U943 : OR2_X1 port map( A1 => mult_143_n6137, A2 => mult_143_n6138, ZN => 
                           n2746);
   U944 : XOR2_X1 port map( A => mult_143_n3455, B => n4657, Z => n2747);
   U948 : XOR2_X1 port map( A => mult_143_n5058, B => mult_143_n5059, Z => 
                           n2755);
   U949 : XOR2_X1 port map( A => mult_143_n4853, B => mult_143_n4852, Z => 
                           n2756);
   U952 : AND2_X1 port map( A1 => n1045, A2 => n1050, ZN => n2757);
   U957 : XOR2_X1 port map( A => mult_143_n4897, B => mult_143_n4896, Z => 
                           n2759);
   U958 : XOR2_X1 port map( A => mult_143_n5067, B => mult_143_n5068, Z => 
                           n2761);
   U959 : OR2_X1 port map( A1 => mult_143_n5532, A2 => mult_143_n5533, ZN => 
                           n2764);
   U961 : AND2_X1 port map( A1 => n3539, A2 => n3789, ZN => n2765);
   U964 : INV_X1 port map( A => mult_143_n812, ZN => mult_143_n6583);
   U965 : AND2_X1 port map( A1 => n671, A2 => n1689, ZN => n2768);
   U966 : INV_X1 port map( A => B_SIG(14), ZN => n865);
   U969 : AND2_X1 port map( A1 => mult_143_n5143, A2 => mult_143_n5144, ZN => 
                           n2769);
   U974 : XOR2_X1 port map( A => A_SIG(11), B => mult_143_n5961, Z => n1744);
   U975 : XNOR2_X1 port map( A => mult_143_n6146, B => mult_143_n6147, ZN => 
                           n1751);
   U976 : XOR2_X1 port map( A => A_SIG(17), B => mult_143_n6012, Z => n1732);
   U983 : OR2_X1 port map( A1 => mult_143_n5132, A2 => mult_143_n5133, ZN => 
                           n1721);
   U987 : XOR2_X1 port map( A => A_SIG(5), B => mult_143_n5862, Z => n1753);
   U988 : XOR2_X1 port map( A => A_SIG(5), B => mult_143_n5860, Z => n1743);
   U989 : XOR2_X1 port map( A => A_SIG(5), B => mult_143_n5864, Z => n1746);
   U992 : XNOR2_X1 port map( A => n4754, B => n1502, ZN => n2778);
   U996 : OR2_X1 port map( A1 => mult_143_n5502, A2 => mult_143_n5503, ZN => 
                           n2784);
   U997 : XOR2_X1 port map( A => mult_143_n5434, B => mult_143_n5435, Z => 
                           n1750);
   U998 : AND2_X1 port map( A1 => mult_143_n5430, A2 => n743, ZN => n2786);
   U1004 : AOI21_X1 port map( B1 => n3756, B2 => n3548, A => n1561, ZN => n2793
                           );
   U1005 : OAI22_X1 port map( A1 => n511, A2 => n512, B1 => mult_143_n5432, B2 
                           => mult_143_n304, ZN => mult_143_n5431);
   U1007 : XNOR2_X1 port map( A => n3605, B => n3730, ZN => n2988);
   U1008 : XNOR2_X1 port map( A => mult_143_n5450, B => n2672, ZN => 
                           mult_143_n5440);
   U1009 : OAI21_X1 port map( B1 => mult_143_n2868, B2 => mult_143_n4493, A => 
                           mult_143_n3154, ZN => mult_143_n393);
   U1011 : XNOR2_X1 port map( A => mult_143_n6040, B => n585, ZN => n1582);
   U1013 : AOI222_X1 port map( A1 => mult_143_n6381, A2 => mult_143_n5419, B1 
                           => mult_143_n6381, B2 => mult_143_n5420, C1 => 
                           mult_143_n5419, C2 => mult_143_n5420, ZN => n2796);
   U1017 : XNOR2_X1 port map( A => mult_143_n5341, B => mult_143_n5338, ZN => 
                           mult_143_n5323);
   U1019 : OAI222_X1 port map( A1 => n4933, A2 => n4581, B1 => n4933, B2 => 
                           n4582, C1 => n4581, C2 => n4582, ZN => n2799);
   U1021 : XNOR2_X1 port map( A => mult_143_n6226, B => n3720, ZN => n2804);
   U1022 : XNOR2_X1 port map( A => n2805, B => n3052, ZN => mult_143_n5592);
   U1023 : XNOR2_X1 port map( A => mult_143_n5905, B => n2864, ZN => n2805);
   U1024 : XOR2_X1 port map( A => mult_143_n5593, B => n711, Z => n2806);
   U1028 : XOR2_X1 port map( A => n2864, B => n2811, Z => mult_143_n1754);
   U1029 : NOR2_X1 port map( A1 => n3644, A2 => n3654, ZN => n2952);
   U1031 : XNOR2_X1 port map( A => mult_143_n5841, B => mult_143_n6367, ZN => 
                           n2812);
   U1032 : INV_X1 port map( A => mult_143_n5048, ZN => n3008);
   U1033 : INV_X1 port map( A => n4622, ZN => n2814);
   U1034 : INV_X1 port map( A => n3064, ZN => n2848);
   U1036 : XNOR2_X1 port map( A => n910, B => mult_143_n6302, ZN => 
                           mult_143_n3094);
   U1039 : XNOR2_X1 port map( A => n2761, B => n2694, ZN => n2970);
   U1044 : XNOR2_X1 port map( A => mult_143_n6040, B => n585, ZN => n1024);
   U1047 : OAI21_X1 port map( B1 => mult_143_n6296, B2 => n909, A => 
                           mult_143_n6308, ZN => n2823);
   U1048 : OAI21_X1 port map( B1 => mult_143_n6296, B2 => n909, A => 
                           mult_143_n6308, ZN => n2824);
   U1049 : NAND2_X1 port map( A1 => n573, A2 => n1077, ZN => n2825);
   U1050 : XNOR2_X1 port map( A => mult_143_n5412, B => mult_143_n5413, ZN => 
                           n1747);
   U1051 : XNOR2_X1 port map( A => n4657, B => mult_143_n5935, ZN => 
                           mult_143_n1724);
   U1053 : XNOR2_X1 port map( A => n2864, B => n2830, ZN => n2829);
   U1055 : NAND2_X1 port map( A1 => mult_143_n5910, A2 => n2955, ZN => n2830);
   U1056 : OAI222_X1 port map( A1 => n2895, A2 => mult_143_n1610, B1 => n4753, 
                           B2 => mult_143_n1553, C1 => mult_143_n1610, C2 => 
                           mult_143_n1553, ZN => n2831);
   U1058 : INV_X1 port map( A => mult_143_n5514, ZN => n3023);
   U1059 : XNOR2_X1 port map( A => n3501, B => n3611, ZN => n1575);
   U1060 : XNOR2_X1 port map( A => mult_143_n5515, B => n3023, ZN => n3022);
   U1064 : AOI222_X1 port map( A1 => n4935, A2 => n3090, B1 => n4935, B2 => 
                           n2730, C1 => n3090, C2 => n2730, ZN => n2835);
   U1065 : AOI222_X1 port map( A1 => n4935, A2 => n3090, B1 => n4935, B2 => 
                           n2730, C1 => n3090, C2 => n2730, ZN => 
                           mult_143_n5554);
   U1068 : XOR2_X1 port map( A => mult_143_n5905, B => n2864, Z => n2837);
   U1071 : XNOR2_X1 port map( A => mult_143_n5987, B => mult_143_n4490, ZN => 
                           n2874);
   U1074 : AOI222_X1 port map( A1 => n969, A2 => n3590, B1 => n969, B2 => 
                           mult_143_n5660, C1 => n3590, C2 => mult_143_n5660, 
                           ZN => mult_143_n5651);
   U1076 : XNOR2_X1 port map( A => n2608, B => mult_143_n6408, ZN => n2844);
   U1078 : NAND2_X1 port map( A1 => n421, A2 => n418, ZN => n2846);
   U1079 : XNOR2_X1 port map( A => n2831, B => n2970, ZN => mult_143_n5468);
   U1081 : OAI222_X1 port map( A1 => n2848, A2 => n2895, B1 => n2848, B2 => 
                           mult_143_n1582, C1 => n4753, C2 => mult_143_n1582, 
                           ZN => n2847);
   U1082 : XNOR2_X1 port map( A => n3018, B => n4632, ZN => n3064);
   U1086 : AOI222_X1 port map( A1 => mult_143_n6382, A2 => n3116, B1 => 
                           mult_143_n6382, B2 => n4607, C1 => n3116, C2 => 
                           n4607, ZN => n2851);
   U1087 : XNOR2_X1 port map( A => n2852, B => mult_143_n5422, ZN => 
                           mult_143_n5166);
   U1088 : XNOR2_X1 port map( A => n2851, B => n961, ZN => n2852);
   U1091 : AND2_X1 port map( A1 => mult_143_n3154, A2 => n4887, ZN => n2855);
   U1093 : INV_X1 port map( A => n740, ZN => n2859);
   U1095 : AOI222_X1 port map( A1 => mult_143_n5511, A2 => mult_143_n5512, B1 
                           => mult_143_n5511, B2 => mult_143_n5510, C1 => 
                           mult_143_n5512, C2 => mult_143_n5510, ZN => n2861);
   U1097 : AOI222_X1 port map( A1 => mult_143_n5511, A2 => mult_143_n5512, B1 
                           => mult_143_n5511, B2 => mult_143_n5510, C1 => 
                           mult_143_n5512, C2 => mult_143_n5510, ZN => 
                           mult_143_n5524);
   U1099 : XNOR2_X1 port map( A => mult_143_n1753, B => n2609, ZN => 
                           mult_143_n5566);
   U1100 : INV_X1 port map( A => n986, ZN => mult_143_n6572);
   U1103 : INV_X1 port map( A => mult_143_n6619, ZN => mult_143_n6496);
   U1106 : XNOR2_X1 port map( A => mult_143_n5974, B => n2895, ZN => n419);
   U1107 : OAI21_X1 port map( B1 => mult_143_n6296, B2 => n909, A => 
                           mult_143_n6308, ZN => mult_143_n6290);
   U1108 : INV_X1 port map( A => mult_143_n1582, ZN => mult_143_n6365);
   U1109 : XNOR2_X1 port map( A => mult_143_n5019, B => n2989, ZN => n3049);
   U1110 : XNOR2_X1 port map( A => mult_143_n5052, B => n2751, ZN => 
                           mult_143_n5048);
   U1115 : NOR2_X1 port map( A1 => n1584, A2 => n3596, ZN => n3021);
   U1123 : OAI22_X1 port map( A1 => mult_143_n5324, A2 => mult_143_n5325, B1 =>
                           mult_143_n5322, B2 => mult_143_n5323, ZN => n2875);
   U1124 : INV_X1 port map( A => mult_143_n1553, ZN => mult_143_n4504);
   U1125 : XNOR2_X1 port map( A => n1683, B => n4829, ZN => n2962);
   U1126 : AOI21_X1 port map( B1 => n2769, B2 => mult_143_n4401, A => n2604, ZN
                           => mult_143_n4788);
   U1127 : XOR2_X1 port map( A => n4657, B => mult_143_n5932, Z => n2877);
   U1129 : XNOR2_X1 port map( A => n4951, B => n1046, ZN => n2881);
   U1133 : XNOR2_X1 port map( A => mult_143_n5950, B => n3803, ZN => n2884);
   U1134 : XNOR2_X1 port map( A => n2812, B => mult_143_n1724, ZN => 
                           mult_143_n5474);
   U1137 : OAI21_X1 port map( B1 => mult_143_n5656, B2 => n3038, A => n3036, ZN
                           => mult_143_n5646);
   U1138 : XNOR2_X1 port map( A => n2679, B => mult_143_n5474, ZN => n2888);
   U1139 : OAI21_X1 port map( B1 => mult_143_n405, B2 => mult_143_n392, A => 
                           mult_143_n393, ZN => n2948);
   U1140 : AOI222_X1 port map( A1 => n3742, A2 => n3510, B1 => n3742, B2 => 
                           n3120, C1 => n3510, C2 => n3120, ZN => n2891);
   U1141 : AOI222_X1 port map( A1 => n3742, A2 => n3510, B1 => n3742, B2 => 
                           n1594, C1 => n1594, C2 => n3510, ZN => mult_143_n430
                           );
   U1142 : NAND4_X1 port map( A1 => n4901, A2 => n2936, A3 => n4936, A4 => 
                           mult_143_n4401, ZN => n618);
   U1144 : XNOR2_X1 port map( A => mult_143_n5592, B => mult_143_n6401, ZN => 
                           n2893);
   U1148 : XNOR2_X1 port map( A => n3097, B => n2895, ZN => mult_143_n1690);
   U1151 : XNOR2_X1 port map( A => n1488, B => n1047, ZN => n2898);
   U1157 : AOI21_X1 port map( B1 => mult_143_n5262, B2 => mult_143_n5261, A => 
                           n386, ZN => n2901);
   U1158 : XNOR2_X1 port map( A => n3556, B => n1839, ZN => mult_143_n4956);
   U1162 : XOR2_X1 port map( A => mult_143_n5479, B => mult_143_n5478, Z => 
                           n2905);
   U1165 : OAI221_X1 port map( B1 => mult_143_n6125, B2 => mult_143_n6126, C1 
                           => mult_143_n6125, C2 => mult_143_n6127, A => 
                           mult_143_n6128, ZN => n2906);
   U1166 : OAI221_X1 port map( B1 => mult_143_n6125, B2 => mult_143_n6126, C1 
                           => mult_143_n6125, C2 => mult_143_n6127, A => 
                           mult_143_n6128, ZN => mult_143_n6036);
   U1167 : INV_X1 port map( A => mult_143_n650, ZN => mult_143_n6581);
   U1168 : NAND2_X1 port map( A1 => n2840, A2 => n3766, ZN => mult_143_n1901);
   U1169 : AND2_X1 port map( A1 => n3775, A2 => n4675, ZN => mult_143_n1528);
   U1170 : XNOR2_X1 port map( A => n3775, B => n3763, ZN => n657);
   U1171 : NAND2_X1 port map( A1 => n3775, A2 => n3827, ZN => n666);
   U1172 : NAND2_X1 port map( A1 => n2600, A2 => mult_143_n5050, ZN => n3009);
   U1178 : AOI21_X1 port map( B1 => n826, B2 => mult_143_n6002, A => 
                           mult_143_n6003, ZN => n2910);
   U1180 : INV_X1 port map( A => mult_143_n4766, ZN => n3002);
   U1183 : XNOR2_X1 port map( A => mult_143_n5669, B => n453, ZN => 
                           mult_143_n5185);
   U1184 : INV_X1 port map( A => n453, ZN => mult_143_n5670);
   U1186 : OAI21_X1 port map( B1 => n632, B2 => n2975, A => n2973, ZN => 
                           mult_143_n6270);
   U1187 : AND2_X1 port map( A1 => mult_143_n6212, A2 => n3044, ZN => 
                           mult_143_n6210);
   U1188 : XOR2_X1 port map( A => mult_143_n5660, B => mult_143_n5661, Z => 
                           n2913);
   U1189 : XNOR2_X1 port map( A => mult_143_n5378, B => n3015, ZN => n3014);
   U1190 : XNOR2_X1 port map( A => n4686, B => n3014, ZN => n1634);
   U1192 : OAI222_X1 port map( A1 => n2770, A2 => n4567, B1 => n4567, B2 => 
                           n2920, C1 => n2770, C2 => n2920, ZN => n2918);
   U1196 : AND2_X1 port map( A1 => mult_143_n5235, A2 => n943, ZN => n2922);
   U1197 : CLKBUF_X1 port map( A => n624, Z => n2923);
   U1198 : AOI22_X1 port map( A1 => n4591, A2 => n4617, B1 => n3809, B2 => 
                           n4714, ZN => n2955);
   U1200 : AOI222_X1 port map( A1 => mult_143_n5651, A2 => mult_143_n5652, B1 
                           => mult_143_n5651, B2 => mult_143_n5650, C1 => 
                           mult_143_n5652, C2 => mult_143_n5650, ZN => n2924);
   U1203 : XNOR2_X1 port map( A => mult_143_n5559, B => n2927, ZN => 
                           mult_143_n5397);
   U1204 : XNOR2_X1 port map( A => mult_143_n5561, B => n4700, ZN => n2927);
   U1217 : AND2_X1 port map( A1 => n3049, A2 => n2675, ZN => n560);
   U1226 : AND2_X1 port map( A1 => n2885, A2 => n821, ZN => n2934);
   U1230 : XNOR2_X1 port map( A => mult_143_n5374, B => n2999, ZN => n2972);
   U1238 : INV_X1 port map( A => n2936, ZN => n956);
   U1239 : XNOR2_X1 port map( A => mult_143_n5483, B => n3034, ZN => n3033);
   U1240 : XNOR2_X1 port map( A => n2937, B => mult_143_n5747, ZN => 
                           mult_143_n5731);
   U1241 : XNOR2_X1 port map( A => n4838, B => n2721, ZN => n2937);
   U1247 : INV_X1 port map( A => mult_143_n5465, ZN => n3041);
   U1248 : XNOR2_X1 port map( A => n2962, B => n3705, ZN => mult_143_n5169);
   U1251 : AOI222_X1 port map( A1 => mult_143_n5181, A2 => mult_143_n5182, B1 
                           => mult_143_n5181, B2 => mult_143_n5180, C1 => 
                           mult_143_n5180, C2 => mult_143_n5182, ZN => n2945);
   U1254 : NAND2_X1 port map( A1 => n4766, A2 => n4665, ZN => n3072);
   U1255 : NAND2_X1 port map( A1 => n3819, A2 => n4766, ZN => n3071);
   U1256 : NAND2_X1 port map( A1 => n3821, A2 => n4765, ZN => n3080);
   U1260 : INV_X1 port map( A => mult_143_n811, ZN => mult_143_n6590);
   U1262 : NAND2_X1 port map( A1 => n4670, A2 => n3768, ZN => mult_143_n5058);
   U1263 : INV_X1 port map( A => n2948, ZN => mult_143_n4767);
   U1264 : XNOR2_X1 port map( A => n4674, B => n3033, ZN => mult_143_n5393);
   U1266 : XNOR2_X1 port map( A => mult_143_n5350, B => n2898, ZN => 
                           mult_143_n5345);
   U1267 : XNOR2_X1 port map( A => n1547, B => n4670, ZN => mult_143_n6479);
   U1268 : NAND2_X1 port map( A1 => n943, A2 => mult_143_n5235, ZN => n963);
   U1269 : AOI21_X1 port map( B1 => mult_143_n4775, B2 => n743, A => n2918, ZN 
                           => mult_143_n4774);
   U1271 : NAND2_X1 port map( A1 => mult_143_n4787, A2 => n824, ZN => n3003);
   U1272 : XNOR2_X1 port map( A => n3769, B => n3579, ZN => mult_143_n6435);
   U1273 : NOR2_X1 port map( A1 => n2951, A2 => n4678, ZN => n441);
   U1275 : NAND2_X1 port map( A1 => n3072, A2 => n2953, ZN => n3018);
   U1282 : NAND2_X1 port map( A1 => n2954, A2 => n1057, ZN => n624);
   U1286 : OAI211_X1 port map( C1 => n3644, C2 => n3657, A => n2957, B => n2956
                           , ZN => mult_143_n5967);
   U1288 : NAND2_X1 port map( A1 => n3778, A2 => n3807, ZN => n2956);
   U1289 : NAND2_X1 port map( A1 => n3777, A2 => n3538, ZN => n2957);
   U1292 : XNOR2_X1 port map( A => n3027, B => n3499, ZN => n1648);
   U1295 : NAND2_X1 port map( A1 => n3003, A2 => n3002, ZN => n720);
   U1297 : AOI21_X1 port map( B1 => n747, B2 => mult_143_n4357, A => 
                           mult_143_n4366, ZN => mult_143_n4771);
   U1298 : NAND2_X1 port map( A1 => mult_143_n4777, A2 => n3004, ZN => 
                           mult_143_n4775);
   U1299 : XNOR2_X1 port map( A => n2960, B => mult_143_n5184, ZN => n1680);
   U1300 : XNOR2_X1 port map( A => mult_143_n5185, B => n4841, ZN => n2960);
   U1302 : NAND2_X1 port map( A1 => n2963, A2 => n2964, ZN => mult_143_n5669);
   U1303 : OR2_X1 port map( A1 => n990, A2 => n4701, ZN => n2963);
   U1305 : NAND2_X1 port map( A1 => n4669, A2 => n4701, ZN => n2964);
   U1309 : INV_X1 port map( A => mult_143_n4401, ZN => n816);
   U1310 : AOI21_X1 port map( B1 => n4578, B2 => n3765, A => n2966, ZN => n1514
                           );
   U1313 : NAND2_X1 port map( A1 => mult_143_n5840, A2 => n2967, ZN => n2966);
   U1314 : NAND2_X1 port map( A1 => n3801, A2 => n3786, ZN => n2967);
   U1319 : INV_X1 port map( A => n666, ZN => mult_143_n1532);
   U1320 : NAND2_X1 port map( A1 => mult_143_n5209, A2 => mult_143_n5208, ZN =>
                           mult_143_n3154);
   U1321 : OAI21_X1 port map( B1 => mult_143_n4828, B2 => mult_143_n2798, A => 
                           n3046, ZN => n3045);
   U1322 : NAND2_X1 port map( A1 => B_SIG(6), A2 => n2978, ZN => n2975);
   U1323 : NAND2_X1 port map( A1 => mult_143_n5071, A2 => n2979, ZN => 
                           mult_143_n5070);
   U1324 : NAND2_X1 port map( A1 => n4672, A2 => n4597, ZN => n2979);
   U1325 : INV_X1 port map( A => mult_143_n686, ZN => mult_143_n6347);
   U1328 : XNOR2_X1 port map( A => mult_143_n5467, B => n3041, ZN => n2980);
   U1330 : NOR2_X1 port map( A1 => mult_143_n5695, A2 => mult_143_n5693, ZN => 
                           n2981);
   U1331 : AOI21_X1 port map( B1 => mult_143_n5695, B2 => mult_143_n5693, A => 
                           n4650, ZN => n2982);
   U1333 : AND2_X1 port map( A1 => n955, A2 => n4657, ZN => n2983);
   U1334 : OAI22_X1 port map( A1 => mult_143_n5699, A2 => n2984, B1 => 
                           mult_143_n5701, B2 => mult_143_n5700, ZN => n1476);
   U1335 : AND2_X1 port map( A1 => mult_143_n5701, A2 => mult_143_n5700, ZN => 
                           n2984);
   U1336 : XNOR2_X1 port map( A => n3603, B => n3490, ZN => n1647);
   U1337 : XNOR2_X1 port map( A => mult_143_n5732, B => mult_143_n5731, ZN => 
                           n2987);
   U1338 : INV_X1 port map( A => mult_143_n5020, ZN => n2989);
   U1339 : NOR2_X1 port map( A1 => n2992, A2 => n2990, ZN => mult_143_n5023);
   U1340 : NAND2_X1 port map( A1 => n595, A2 => n2991, ZN => n2990);
   U1341 : NAND2_X1 port map( A1 => n4589, A2 => n3641, ZN => n2991);
   U1342 : INV_X1 port map( A => mult_143_n5025, ZN => n2992);
   U1343 : NOR2_X1 port map( A1 => n2803, A2 => mult_143_n6432, ZN => n2993);
   U1344 : XNOR2_X1 port map( A => mult_143_n5252, B => n2995, ZN => n1570);
   U1345 : XNOR2_X1 port map( A => mult_143_n5250, B => n2996, ZN => n2995);
   U1346 : INV_X1 port map( A => mult_143_n5251, ZN => n2996);
   U1347 : NAND2_X1 port map( A1 => n2901, A2 => n2997, ZN => mult_143_n5257);
   U1348 : AND2_X1 port map( A1 => mult_143_n5266, A2 => mult_143_n5265, ZN => 
                           n2997);
   U1350 : NAND2_X1 port map( A1 => mult_143_n4954, A2 => n2998, ZN => 
                           mult_143_n4953);
   U1351 : NAND2_X1 port map( A1 => n4672, A2 => n4576, ZN => n2998);
   U1352 : INV_X1 port map( A => mult_143_n5375, ZN => n2999);
   U1353 : XNOR2_X1 port map( A => mult_143_n5893, B => n3099, ZN => 
                           mult_143_n6421);
   U1354 : AND2_X1 port map( A1 => n1590, A2 => n1614, ZN => n3001);
   U1355 : INV_X1 port map( A => n720, ZN => mult_143_n4784);
   U1356 : OAI21_X1 port map( B1 => n3535, B2 => n3813, A => n4612, ZN => n1541
                           );
   U1357 : OR2_X1 port map( A1 => mult_143_n5050, A2 => n2600, ZN => n3006);
   U1358 : NAND2_X1 port map( A1 => n3009, A2 => n3008, ZN => n3007);
   U1359 : XNOR2_X1 port map( A => n3600, B => n3593, ZN => n1678);
   U1360 : XNOR2_X1 port map( A => mult_143_n5401, B => n4758, ZN => n3010);
   U1361 : NAND2_X1 port map( A1 => n3012, A2 => n3011, ZN => mult_143_n5387);
   U1362 : OR2_X1 port map( A1 => n3013, A2 => mult_143_n5389, ZN => n3011);
   U1363 : NAND2_X1 port map( A1 => mult_143_n5389, A2 => n3013, ZN => n3012);
   U1364 : INV_X1 port map( A => n966, ZN => n3013);
   U1365 : INV_X1 port map( A => mult_143_n5377, ZN => n3015);
   U1367 : XNOR2_X1 port map( A => mult_143_n5724, B => n3017, ZN => n3016);
   U1368 : INV_X1 port map( A => mult_143_n5723, ZN => n3017);
   U1369 : XNOR2_X1 port map( A => mult_143_n6435, B => n3019, ZN => 
                           mult_143_n5347);
   U1370 : XNOR2_X1 port map( A => n2689, B => n1752, ZN => n3019);
   U1372 : NOR2_X1 port map( A1 => n2722, A2 => n3021, ZN => n3020);
   U1373 : NAND2_X1 port map( A1 => mult_143_n5765, A2 => n3025, ZN => n3024);
   U1374 : NAND2_X1 port map( A1 => mult_143_n6347, A2 => mult_143_n6348, ZN =>
                           n3025);
   U1376 : XNOR2_X1 port map( A => mult_143_n5653, B => n2913, ZN => n3026);
   U1377 : INV_X1 port map( A => mult_143_n5019, ZN => n3029);
   U1378 : OAI21_X1 port map( B1 => n4857, B2 => n3032, A => n3031, ZN => 
                           mult_143_n5702);
   U1379 : OR2_X1 port map( A1 => mult_143_n5689, A2 => mult_143_n5690, ZN => 
                           n3031);
   U1380 : AND2_X1 port map( A1 => mult_143_n5689, A2 => mult_143_n5690, ZN => 
                           n3032);
   U1381 : INV_X1 port map( A => mult_143_n5481, ZN => n3034);
   U1382 : OAI211_X1 port map( C1 => n3527, C2 => n3554, A => n3668, B => n3601
                           , ZN => n1520);
   U1384 : NAND2_X1 port map( A1 => n3037, A2 => mult_143_n812, ZN => n3036);
   U1385 : INV_X1 port map( A => mult_143_n5658, ZN => n3037);
   U1386 : AND2_X1 port map( A1 => mult_143_n5658, A2 => mult_143_n6583, ZN => 
                           n3038);
   U1387 : NOR2_X1 port map( A1 => mult_143_n5058, A2 => n3824, ZN => n3039);
   U1388 : XNOR2_X1 port map( A => mult_143_n4490, B => n4603, ZN => n3042);
   U1390 : INV_X1 port map( A => n3045, ZN => n3044);
   U1391 : NAND2_X1 port map( A1 => mult_143_n48, A2 => B_SIG(5), ZN => n3046);
   U1394 : INV_X1 port map( A => n955, ZN => mult_143_n6605);
   U1397 : XNOR2_X1 port map( A => mult_143_n5854, B => n3791, ZN => n3052);
   U1398 : AND2_X1 port map( A1 => n3079, A2 => n3080, ZN => n3053);
   U1399 : XNOR2_X1 port map( A => n4750, B => mult_143_n6066, ZN => n3054);
   U1400 : AND2_X1 port map( A1 => n3077, A2 => n3078, ZN => n3055);
   U1401 : XNOR2_X1 port map( A => n4750, B => mult_143_n6067, ZN => n3056);
   U1402 : XNOR2_X1 port map( A => mult_143_n5855, B => n3791, ZN => n3057);
   U1403 : XOR2_X1 port map( A => mult_143_n4490, B => mult_143_n6008, Z => 
                           n3058);
   U1404 : XNOR2_X1 port map( A => mult_143_n5959, B => n3793, ZN => n3059);
   U1405 : AND2_X1 port map( A1 => n3075, A2 => n3076, ZN => n3060);
   U1406 : XOR2_X1 port map( A => mult_143_n1891, B => n4750, Z => n3061);
   U1407 : NAND2_X1 port map( A1 => n2840, A2 => n4766, ZN => mult_143_n1891);
   U1408 : XNOR2_X1 port map( A => mult_143_n5914, B => n3792, ZN => n3062);
   U1409 : AND2_X1 port map( A1 => n3073, A2 => n3074, ZN => n3063);
   U1410 : XNOR2_X1 port map( A => n4760, B => mult_143_n6047, ZN => n3065);
   U1412 : XNOR2_X1 port map( A => mult_143_n5986, B => n3794, ZN => n3067);
   U1413 : AND2_X1 port map( A1 => n3069, A2 => n3070, ZN => n3068);
   U1415 : NOR2_X1 port map( A1 => n2633, A2 => n2751, ZN => mult_143_n5778);
   U1416 : INV_X1 port map( A => mult_143_n1892, ZN => mult_143_n1521);
   U1417 : INV_X1 port map( A => mult_143_n1894, ZN => mult_143_n1523);
   U1418 : INV_X1 port map( A => mult_143_n1901, ZN => mult_143_n1530);
   U1419 : NAND2_X1 port map( A1 => n3820, A2 => n4766, ZN => n3070);
   U1420 : NAND2_X1 port map( A1 => n2814, A2 => n3804, ZN => n3069);
   U1421 : NAND2_X1 port map( A1 => n3798, A2 => n4766, ZN => mult_143_n2200);
   U1422 : NAND2_X1 port map( A1 => n3533, A2 => n4766, ZN => mult_143_n2066);
   U1423 : NAND2_X1 port map( A1 => n2840, A2 => n4890, ZN => mult_143_n1897);
   U1424 : NAND2_X1 port map( A1 => n3775, A2 => n3804, ZN => mult_143_n1892);
   U1425 : NAND2_X1 port map( A1 => n3809, A2 => n4766, ZN => n3074);
   U1426 : NAND2_X1 port map( A1 => n3536, A2 => n3804, ZN => n3073);
   U1427 : NAND2_X1 port map( A1 => n3817, A2 => n4766, ZN => n3076);
   U1428 : NAND2_X1 port map( A1 => n3799, A2 => n3804, ZN => n3075);
   U1429 : NAND2_X1 port map( A1 => n3799, A2 => n4766, ZN => mult_143_n2267);
   U1430 : NAND2_X1 port map( A1 => n3539, A2 => n4766, ZN => mult_143_n2133);
   U1431 : NAND2_X1 port map( A1 => n3771, A2 => n4766, ZN => mult_143_n2401);
   U1432 : NAND2_X1 port map( A1 => n3540, A2 => n4766, ZN => mult_143_n2001);
   U1433 : NAND2_X1 port map( A1 => n3806, A2 => n4765, ZN => n3078);
   U1434 : NAND2_X1 port map( A1 => n3540, A2 => n3804, ZN => n3077);
   U1435 : NAND2_X1 port map( A1 => n3771, A2 => n3789, ZN => n3079);
   U1436 : NAND2_X1 port map( A1 => n2840, A2 => n4695, ZN => mult_143_n1896);
   U1437 : NAND2_X1 port map( A1 => n2840, A2 => n2908, ZN => mult_143_n1894);
   U1438 : NAND2_X1 port map( A1 => n2840, A2 => n4871, ZN => mult_143_n1893);
   U21 : BUF_X1 port map( A => mult_143_n4755, Z => n2947);
   U187 : XOR2_X1 port map( A => A_SIG(3), B => A_SIG(2), Z => mult_143_n6199);
   U430 : XNOR2_X1 port map( A => A_SIG(3), B => A_SIG(4), ZN => mult_143_n6200
                           );
   U226 : NAND2_X1 port map( A1 => B_SIG(13), A2 => B_SIG(11), ZN => n2971);
   mult_143_U4659 : XOR2_X1 port map( A => A_SIG(6), B => A_SIG(5), Z => 
                           mult_143_n6254);
   U770 : NAND2_X1 port map( A1 => mult_143_n6199, A2 => mult_143_n6198, ZN => 
                           mult_143_n5859);
   U728 : NAND2_X1 port map( A1 => n650, A2 => mult_143_n6306, ZN => 
                           mult_143_n4824);
   U1395 : OR2_X1 port map( A1 => n2751, A2 => n3051, ZN => n3050);
   U973 : INV_X1 port map( A => B_SIG(13), ZN => n868);
   U361 : INV_X1 port map( A => A_SIG(11), ZN => n1765);
   U505 : INV_X1 port map( A => B_SIG(11), ZN => n874);
   mult_143_U4021 : AND3_X1 port map( A1 => mult_143_n6306, A2 => 
                           mult_143_n6305, A3 => mult_143_n6231, ZN => 
                           mult_143_n72);
   U1332 : NOR2_X1 port map( A1 => mult_143_n5712, A2 => n2983, ZN => 
                           mult_143_n5695);
   U44 : NAND2_X1 port map( A1 => n3083, A2 => n3082, ZN => mult_143_n5394);
   U54 : OR2_X1 port map( A1 => mult_143_n5374, A2 => mult_143_n5375, ZN => 
                           n3082);
   U59 : NAND2_X1 port map( A1 => n3084, A2 => n3085, ZN => n3083);
   U79 : INV_X1 port map( A => mult_143_n5372, ZN => n3085);
   U83 : OAI211_X1 port map( C1 => n3613, C2 => n3659, A => n3087, B => n3086, 
                           ZN => mult_143_n5842);
   U84 : NAND2_X1 port map( A1 => n3786, A2 => n3821, ZN => n3086);
   U87 : NAND2_X1 port map( A1 => n4695, A2 => n3771, ZN => n3087);
   U148 : AOI222_X1 port map( A1 => n2806, A2 => n2893, B1 => mult_143_n5570, 
                           B2 => n2806, C1 => mult_143_n5570, C2 => n2893, ZN 
                           => mult_143_n5574);
   U184 : AOI222_X1 port map( A1 => n962, A2 => mult_143_n5381, B1 => n962, B2 
                           => mult_143_n5380, C1 => mult_143_n5381, C2 => 
                           mult_143_n5380, ZN => mult_143_n5378);
   U288 : NAND2_X1 port map( A1 => mult_143_n5828, A2 => n3122, ZN => n3121);
   U336 : INV_X1 port map( A => n997, ZN => n2598);
   U344 : NOR2_X1 port map( A1 => mult_143_n5945, A2 => n3129, ZN => 
                           mult_143_n5944);
   U349 : NOR2_X1 port map( A1 => mult_143_n5936, A2 => n2958, ZN => 
                           mult_143_n5935);
   U369 : OR2_X1 port map( A1 => n648, A2 => mult_143_n6292, ZN => n979);
   U454 : AND2_X1 port map( A1 => n4890, A2 => n3817, ZN => n3129);
   U476 : XNOR2_X1 port map( A => n3740, B => n4592, ZN => n3135);
   U483 : NOR2_X1 port map( A1 => mult_143_n6092, A2 => n3132, ZN => n3131);
   U488 : XNOR2_X1 port map( A => mult_143_n6216, B => n3135, ZN => n1047);
   U509 : OAI21_X1 port map( B1 => B_SIG(11), B2 => B_SIG(13), A => B_SIG(12), 
                           ZN => n1072);
   U597 : XNOR2_X1 port map( A => n3131, B => n4752, ZN => n2732);
   U699 : INV_X1 port map( A => B_SIG(4), ZN => n2977);
   U807 : NAND2_X1 port map( A1 => mult_143_n5813, A2 => n3126, ZN => n3125);
   U883 : XNOR2_X1 port map( A => mult_143_n5505, B => n3134, ZN => n3133);
   U891 : XOR2_X1 port map( A => A_SIG(4), B => A_SIG(5), Z => mult_143_n6198);
   U921 : XNOR2_X1 port map( A => A_SIG(17), B => A_SIG(18), ZN => 
                           mult_143_n6293);
   U947 : AOI21_X1 port map( B1 => n3127, B2 => n3123, A => n3125, ZN => 
                           mult_143_n5811);
   U994 : OAI22_X1 port map( A1 => mult_143_n5683, A2 => n3128, B1 => 
                           mult_143_n5686, B2 => mult_143_n5685, ZN => 
                           mult_143_n5699);
   U1052 : AOI222_X1 port map( A1 => n3115, A2 => n975, B1 => n3115, B2 => 
                           mult_143_n5786, C1 => n975, C2 => mult_143_n5786, ZN
                           => mult_143_n5776);
   U1054 : XOR2_X1 port map( A => A_SIG(17), B => A_SIG(16), Z => 
                           mult_143_n6306);
   U1069 : INV_X1 port map( A => A_SIG(2), ZN => n536);
   U1070 : AND3_X1 port map( A1 => mult_143_n6110, A2 => mult_143_n4832, A3 => 
                           mult_143_n6111, ZN => mult_143_n96);
   U1077 : AOI21_X1 port map( B1 => n4620, B2 => n3765, A => n3121, ZN => n1537
                           );
   U1080 : NAND2_X1 port map( A1 => n648, A2 => mult_143_n6284, ZN => 
                           mult_143_n4820);
   U1098 : INV_X1 port map( A => mult_143_n5647, ZN => n3138);
   U1149 : AOI22_X1 port map( A1 => n986, A2 => n1657, B1 => n496, B2 => n1042,
                           ZN => n3093);
   U1150 : AOI21_X1 port map( B1 => mult_143_n6022, B2 => mult_143_n6030, A => 
                           mult_143_n6031, ZN => n3095);
   U1176 : XNOR2_X1 port map( A => mult_143_n5048, B => n3100, ZN => n2613);
   U1202 : XNOR2_X1 port map( A => mult_143_n5050, B => n2600, ZN => n3100);
   U1231 : INV_X1 port map( A => A_SIG(5), ZN => n642);
   U1234 : AOI222_X1 port map( A1 => n2715, A2 => n4839, B1 => n2715, B2 => 
                           mult_143_n5463, C1 => n4839, C2 => mult_143_n5463, 
                           ZN => n3101);
   U1246 : XNOR2_X1 port map( A => mult_143_n5569, B => mult_143_n5570, ZN => 
                           n3104);
   U1258 : AOI21_X1 port map( B1 => mult_143_n6022, B2 => mult_143_n6030, A => 
                           mult_143_n6031, ZN => mult_143_n5939);
   U1265 : XOR2_X1 port map( A => n4658, B => n608, Z => n3105);
   U1283 : XOR2_X1 port map( A => n4658, B => n608, Z => n3106);
   U1308 : XOR2_X1 port map( A => mult_143_n5971, B => n2895, Z => n3107);
   U1315 : AOI222_X1 port map( A1 => n4658, A2 => n4630, B1 => n4658, B2 => 
                           mult_143_n4937, C1 => mult_143_n4937, C2 => n4630, 
                           ZN => n3108);
   U1329 : AOI222_X1 port map( A1 => n4658, A2 => n4630, B1 => mult_143_n4939, 
                           B2 => mult_143_n4937, C1 => mult_143_n4937, C2 => 
                           n4630, ZN => n990);
   U1414 : XNOR2_X1 port map( A => n4856, B => mult_143_n5600, ZN => 
                           mult_143_n5588);
   U1440 : XNOR2_X1 port map( A => n617, B => n1049, ZN => n3110);
   U1443 : XOR2_X1 port map( A => n4657, B => mult_143_n5935, Z => n3112);
   U1446 : AOI222_X1 port map( A1 => n2726, A2 => n3795, B1 => n2726, B2 => 
                           n3050, C1 => n3795, C2 => n3050, ZN => n3115);
   U1454 : NAND2_X1 port map( A1 => n3801, A2 => n4675, ZN => n3122);
   U1455 : INV_X1 port map( A => mult_143_n5124, ZN => n3123);
   U1456 : NAND2_X1 port map( A1 => mult_143_n2, A2 => B_SIG(10), ZN => n3126);
   U1457 : INV_X1 port map( A => mult_143_n6627, ZN => n3127);
   U1458 : AND2_X1 port map( A1 => mult_143_n5685, A2 => mult_143_n5686, ZN => 
                           n3128);
   U1459 : OR2_X1 port map( A1 => mult_143_n2702, A2 => mult_143_n1719, ZN => 
                           mult_143_n5621);
   U1460 : AND2_X1 port map( A1 => n1624, A2 => n1625, ZN => n3130);
   U1461 : AND2_X1 port map( A1 => n2908, A2 => n3820, ZN => n3132);
   U1462 : XNOR2_X1 port map( A => n3133, B => mult_143_n5507, ZN => n1638);
   U1463 : INV_X1 port map( A => mult_143_n5508, ZN => n3134);
   U1464 : AND2_X1 port map( A1 => mult_143_n1690, A2 => mult_143_n1754, ZN => 
                           mult_143_n5591);
   U1465 : OAI211_X1 port map( C1 => n3644, C2 => n3665, A => n3137, B => n3136
                           , ZN => mult_143_n5972);
   U1466 : NAND2_X1 port map( A1 => n3779, A2 => n3807, ZN => n3136);
   U1467 : NAND2_X1 port map( A1 => n3827, A2 => n3538, ZN => n3137);
   U1468 : NOR2_X1 port map( A1 => mult_143_n5912, A2 => n3140, ZN => n3139);
   U1469 : AND2_X1 port map( A1 => n3804, A2 => n3809, ZN => n3140);
   U1470 : OAI211_X1 port map( C1 => mult_143_n4842, C2 => mult_143_n3443, A =>
                           n3142, B => n3141, ZN => mult_143_n4963);
   U1471 : NAND2_X1 port map( A1 => B_SIG(14), A2 => mult_143_n74, ZN => n3141)
                           ;
   U1472 : NAND2_X1 port map( A1 => B_SIG(12), A2 => mult_143_n84, ZN => n3142)
                           ;
   U1473 : OAI21_X1 port map( B1 => n3143, B2 => mult_143_n4766, A => n1038, ZN
                           => n2954);
   U1474 : AOI21_X1 port map( B1 => n620, B2 => mult_143_n4767, A => n618, ZN 
                           => n3143);
   MY_CLK_r_REG1510_S1 : DFF_X1 port map( D => n1724, CK => clk, Q => n3831, QN
                           => n_1170);
   MY_CLK_r_REG1164_S2 : DFF_X1 port map( D => n1836, CK => clk, Q => n3830, QN
                           => n_1171);
   MY_CLK_r_REG1262_S2 : DFF_X1 port map( D => n718, CK => clk, Q => n3829, QN 
                           => n4855);
   MY_CLK_r_REG1125_S3 : DFF_X1 port map( D => n747, CK => clk, Q => n3828, QN 
                           => n_1172);
   MY_CLK_r_REG1253_S1 : DFF_X1 port map( D => n1832, CK => clk, Q => n3826, QN
                           => n4624);
   MY_CLK_r_REG1343_S1 : DFF_X1 port map( D => n772, CK => clk, Q => n3825, QN 
                           => n_1173);
   MY_CLK_r_REG1509_S1 : DFF_X1 port map( D => n1828, CK => clk, Q => n3824, QN
                           => n4603);
   MY_CLK_r_REG1416_S1 : DFF_X1 port map( D => n755, CK => clk, Q => n3823, QN 
                           => n_1174);
   MY_CLK_r_REG1503_S1 : DFF_X1 port map( D => n688, CK => clk, Q => n3822, QN 
                           => n_1175);
   MY_CLK_r_REG1470_S1 : DFF_X1 port map( D => mult_143_n3245, CK => clk, Q => 
                           n3821, QN => n_1176);
   MY_CLK_r_REG1297_S1 : DFF_X1 port map( D => n799, CK => clk, Q => n3820, QN 
                           => n_1177);
   MY_CLK_r_REG1355_S1 : DFF_X1 port map( D => n774, CK => clk, Q => n3819, QN 
                           => n_1178);
   MY_CLK_r_REG1185_S2 : DFF_X1 port map( D => n1787, CK => clk, Q => n3818, QN
                           => n_1179);
   MY_CLK_r_REG1427_S1 : DFF_X1 port map( D => n1023, CK => clk, Q => n3817, QN
                           => n_1180);
   MY_CLK_r_REG1261_S1 : DFF_X1 port map( D => n1722, CK => clk, Q => n3816, QN
                           => n_1181);
   MY_CLK_r_REG1251_S1 : DFF_X1 port map( D => n1723, CK => clk, Q => n3815, QN
                           => n_1182);
   MY_CLK_r_REG1252_S1 : DFF_X1 port map( D => n1728, CK => clk, Q => n3814, QN
                           => n_1183);
   MY_CLK_r_REG1209_S3 : DFF_X1 port map( D => mult_143_n6535, CK => clk, Q => 
                           n3813, QN => n_1184);
   MY_CLK_r_REG1240_S3 : DFF_X1 port map( D => mult_143_n6524, CK => clk, Q => 
                           n3812, QN => n_1185);
   MY_CLK_r_REG1428_S1 : DFF_X1 port map( D => n1759, CK => clk, Q => n3811, QN
                           => n_1186);
   MY_CLK_r_REG1319_S1 : DFF_X1 port map( D => n778, CK => clk, Q => n3810, QN 
                           => n4738);
   MY_CLK_r_REG1452_S1 : DFF_X1 port map( D => n1031, CK => clk, Q => n3809, QN
                           => n_1187);
   MY_CLK_r_REG1402_S1 : DFF_X1 port map( D => n787, CK => clk, Q => n3807, QN 
                           => n4629);
   MY_CLK_r_REG1326_S1 : DFF_X1 port map( D => n1027, CK => clk, Q => n3806, QN
                           => n_1188);
   MY_CLK_r_REG1465_S1 : DFF_X1 port map( D => mult_143_n2, CK => clk, Q => 
                           n3801, QN => n_1189);
   MY_CLK_r_REG1425_S1 : DFF_X1 port map( D => mult_143_n36, CK => clk, Q => 
                           n3799, QN => n_1190);
   MY_CLK_r_REG1400_S1 : DFF_X1 port map( D => mult_143_n48, CK => clk, Q => 
                           n3798, QN => n_1191);
   MY_CLK_r_REG1358_S1 : DFF_X1 port map( D => A_SIG(14), CK => clk, Q => n3795
                           , QN => n4634);
   MY_CLK_r_REG1405_S1 : DFF_X1 port map( D => A_SIG(8), CK => clk, Q => n3793,
                           QN => n4625);
   MY_CLK_r_REG1453_S1 : DFF_X1 port map( D => A_SIG(2), CK => clk, Q => n3791,
                           QN => n4630);
   MY_CLK_r_REG1496_S1 : DFF_X1 port map( D => B_SIG(13), CK => clk, Q => n3780
                           , QN => n_1192);
   MY_CLK_r_REG1506_S1 : DFF_X1 port map( D => B_SIG(10), CK => clk, Q => n3778
                           , QN => n_1193);
   MY_CLK_r_REG1507_S1 : DFF_X1 port map( D => B_SIG(9), CK => clk, Q => n3777,
                           QN => n_1194);
   MY_CLK_r_REG1499_S1 : DFF_X1 port map( D => B_SIG(13), CK => clk, Q => n3766
                           , QN => n_1195);
   MY_CLK_r_REG1463_S1 : DFF_X1 port map( D => n3123, CK => clk, Q => n3765, QN
                           => n_1196);
   MY_CLK_r_REG1382_S1 : DFF_X1 port map( D => n4623, CK => clk, Q => n3764, QN
                           => n_1197);
   MY_CLK_r_REG1192_S1 : DFF_X1 port map( D => n2706, CK => clk, Q => n3763, QN
                           => n_1198);
   MY_CLK_r_REG1469_S1 : DFF_X1 port map( D => mult_143_n3245, CK => clk, Q => 
                           n3762, QN => n_1199);
   MY_CLK_r_REG1434_S1 : DFF_X1 port map( D => n1715, CK => clk, Q => n3761, QN
                           => n_1200);
   MY_CLK_r_REG1430_S1 : DFF_X1 port map( D => n1713, CK => clk, Q => n3759, QN
                           => n4618);
   MY_CLK_r_REG1245_S2 : DFF_X1 port map( D => mult_143_n5789, CK => clk, Q => 
                           n3758, QN => n_1201);
   MY_CLK_r_REG1243_S2 : DFF_X1 port map( D => mult_143_n5788, CK => clk, Q => 
                           n3757, QN => n_1202);
   MY_CLK_r_REG1298_S1 : DFF_X1 port map( D => mult_143_n994, CK => clk, Q => 
                           n_1203, QN => n4575);
   MY_CLK_r_REG1195_S2 : DFF_X1 port map( D => n1708, CK => clk, Q => n3754, QN
                           => n_1204);
   MY_CLK_r_REG1191_S2 : DFF_X1 port map( D => mult_143_n5158, CK => clk, Q => 
                           n_1205, QN => n4826);
   MY_CLK_r_REG1163_S2 : DFF_X1 port map( D => n1707, CK => clk, Q => n3752, QN
                           => n_1206);
   MY_CLK_r_REG1236_S2 : DFF_X1 port map( D => n1706, CK => clk, Q => n3751, QN
                           => n_1207);
   MY_CLK_r_REG1220_S2 : DFF_X1 port map( D => n1705, CK => clk, Q => n3750, QN
                           => n_1208);
   MY_CLK_r_REG1145_S2 : DFF_X1 port map( D => mult_143_n5576, CK => clk, Q => 
                           n3749, QN => n4903);
   MY_CLK_r_REG1365_S1 : DFF_X1 port map( D => n1703, CK => clk, Q => n3748, QN
                           => n_1209);
   MY_CLK_r_REG1221_S2 : DFF_X1 port map( D => n1701, CK => clk, Q => n3746, QN
                           => n4639);
   MY_CLK_r_REG1172_S2 : DFF_X1 port map( D => n1700, CK => clk, Q => n3745, QN
                           => n_1210);
   MY_CLK_r_REG1223_S3 : DFF_X1 port map( D => mult_143_n4756, CK => clk, Q => 
                           n3744, QN => n_1211);
   MY_CLK_r_REG1208_S3 : DFF_X1 port map( D => mult_143_n4773, CK => clk, Q => 
                           n3743, QN => n_1212);
   MY_CLK_r_REG1372_S1 : DFF_X1 port map( D => mult_143_n6201, CK => clk, Q => 
                           n3741, QN => n_1213);
   MY_CLK_r_REG1366_S1 : DFF_X1 port map( D => n1695, CK => clk, Q => n3740, QN
                           => n_1214);
   MY_CLK_r_REG1143_S2 : DFF_X1 port map( D => mult_143_n5216, CK => clk, Q => 
                           n3739, QN => n_1215);
   MY_CLK_r_REG1231_S2 : DFF_X1 port map( D => n1688, CK => clk, Q => n3737, QN
                           => n4725);
   MY_CLK_r_REG1235_S2 : DFF_X1 port map( D => mult_143_n5698, CK => clk, Q => 
                           n3736, QN => n_1216);
   MY_CLK_r_REG1183_S2 : DFF_X1 port map( D => n1686, CK => clk, Q => n3735, QN
                           => n_1217);
   MY_CLK_r_REG1178_S2 : DFF_X1 port map( D => n1685, CK => clk, Q => n3734, QN
                           => n_1218);
   MY_CLK_r_REG1257_S2 : DFF_X1 port map( D => mult_143_n5679, CK => clk, Q => 
                           n3732, QN => n4852);
   MY_CLK_r_REG1196_S2 : DFF_X1 port map( D => mult_143_n5159, CK => clk, Q => 
                           n3731, QN => n_1219);
   MY_CLK_r_REG1188_S2 : DFF_X1 port map( D => n1681, CK => clk, Q => n3730, QN
                           => n_1220);
   MY_CLK_r_REG1367_S1 : DFF_X1 port map( D => n1679, CK => clk, Q => n3729, QN
                           => n_1221);
   MY_CLK_r_REG1205_S2 : DFF_X1 port map( D => n1676, CK => clk, Q => n3728, QN
                           => n4869);
   MY_CLK_r_REG1204_S2 : DFF_X1 port map( D => mult_143_n5613, CK => clk, Q => 
                           n_1222, QN => n4849);
   MY_CLK_r_REG1371_S1 : DFF_X1 port map( D => mult_143_n6264, CK => clk, Q => 
                           n3725, QN => n_1223);
   MY_CLK_r_REG1194_S1 : DFF_X1 port map( D => n1674, CK => clk, Q => n3724, QN
                           => n4599);
   MY_CLK_r_REG1333_S1 : DFF_X1 port map( D => n1672, CK => clk, Q => n3723, QN
                           => n_1224);
   MY_CLK_r_REG1340_S1 : DFF_X1 port map( D => mult_143_n6263, CK => clk, Q => 
                           n3722, QN => n_1225);
   MY_CLK_r_REG1339_S1 : DFF_X1 port map( D => n1668, CK => clk, Q => n3721, QN
                           => n_1226);
   MY_CLK_r_REG1338_S1 : DFF_X1 port map( D => n1667, CK => clk, Q => n3720, QN
                           => n_1227);
   MY_CLK_r_REG1389_S1 : DFF_X1 port map( D => n1666, CK => clk, Q => n3719, QN
                           => n4592);
   MY_CLK_r_REG1388_S1 : DFF_X1 port map( D => mult_143_n6203, CK => clk, Q => 
                           n3718, QN => n_1228);
   MY_CLK_r_REG1413_S1 : DFF_X1 port map( D => n1663, CK => clk, Q => n3717, QN
                           => n4581);
   MY_CLK_r_REG1387_S1 : DFF_X1 port map( D => n1662, CK => clk, Q => n3716, QN
                           => n4582);
   MY_CLK_r_REG1359_S1 : DFF_X1 port map( D => mult_143_n6168, CK => clk, Q => 
                           n3715, QN => n_1229);
   MY_CLK_r_REG1386_S1 : DFF_X1 port map( D => n1661, CK => clk, Q => n3714, QN
                           => n4627);
   MY_CLK_r_REG1412_S1 : DFF_X1 port map( D => n1660, CK => clk, Q => n3713, QN
                           => n4655);
   MY_CLK_r_REG1381_S1 : DFF_X1 port map( D => n1659, CK => clk, Q => n3712, QN
                           => n4584);
   MY_CLK_r_REG1218_S2 : DFF_X1 port map( D => n1650, CK => clk, Q => n3711, QN
                           => n_1230);
   MY_CLK_r_REG1230_S2 : DFF_X1 port map( D => mult_143_n5466, CK => clk, Q => 
                           n_1231, QN => n4964);
   MY_CLK_r_REG1224_S2 : DFF_X1 port map( D => n1649, CK => clk, Q => n3709, QN
                           => n_1232);
   MY_CLK_r_REG1225_S2 : DFF_X1 port map( D => n1646, CK => clk, Q => n3707, QN
                           => n_1233);
   MY_CLK_r_REG1166_S2 : DFF_X1 port map( D => n1643, CK => clk, Q => n3705, QN
                           => n4636);
   MY_CLK_r_REG1200_S2 : DFF_X1 port map( D => mult_143_n5620, CK => clk, Q => 
                           n_1234, QN => n4850);
   MY_CLK_r_REG1147_S2 : DFF_X1 port map( D => mult_143_n5614, CK => clk, Q => 
                           n3703, QN => n_1235);
   MY_CLK_r_REG1198_S2 : DFF_X1 port map( D => mult_143_n5215, CK => clk, Q => 
                           n3702, QN => n4895);
   MY_CLK_r_REG1242_S2 : DFF_X1 port map( D => n1640, CK => clk, Q => n3700, QN
                           => n_1236);
   MY_CLK_r_REG1241_S2 : DFF_X1 port map( D => n1639, CK => clk, Q => n3699, QN
                           => n4637);
   MY_CLK_r_REG1337_S1 : DFF_X1 port map( D => n1637, CK => clk, Q => n3698, QN
                           => n_1237);
   MY_CLK_r_REG1311_S1 : DFF_X1 port map( D => n1636, CK => clk, Q => n3697, QN
                           => n4702);
   MY_CLK_r_REG1207_S2 : DFF_X1 port map( D => n1635, CK => clk, Q => n3696, QN
                           => n_1238);
   MY_CLK_r_REG1206_S1 : DFF_X1 port map( D => mult_143_n4850, CK => clk, Q => 
                           n3695, QN => n_1239);
   MY_CLK_r_REG1457_S1 : DFF_X1 port map( D => mult_143_n5117, CK => clk, Q => 
                           n3694, QN => n_1240);
   MY_CLK_r_REG1431_S1 : DFF_X1 port map( D => mult_143_n5118, CK => clk, Q => 
                           n3693, QN => n_1241);
   MY_CLK_r_REG1406_S1 : DFF_X1 port map( D => n1630, CK => clk, Q => n3692, QN
                           => n4601);
   MY_CLK_r_REG1202_S1 : DFF_X1 port map( D => n1622, CK => clk, Q => n3691, QN
                           => n_1242);
   MY_CLK_r_REG1407_S1 : DFF_X1 port map( D => n1618, CK => clk, Q => n3690, QN
                           => n_1243);
   MY_CLK_r_REG1336_S1 : DFF_X1 port map( D => n1616, CK => clk, Q => n3689, QN
                           => n_1244);
   MY_CLK_r_REG1415_S1 : DFF_X1 port map( D => mult_143_n5318, CK => clk, Q => 
                           n3688, QN => n_1245);
   MY_CLK_r_REG1483_S1 : DFF_X1 port map( D => n1557, CK => clk, Q => n3687, QN
                           => n4626);
   MY_CLK_r_REG1327_S1 : DFF_X1 port map( D => n1612, CK => clk, Q => n3686, QN
                           => n_1246);
   MY_CLK_r_REG1356_S1 : DFF_X1 port map( D => n1611, CK => clk, Q => n3685, QN
                           => n4610);
   MY_CLK_r_REG1433_S1 : DFF_X1 port map( D => n1609, CK => clk, Q => n3683, QN
                           => n4613);
   MY_CLK_r_REG1309_S1 : DFF_X1 port map( D => n1608, CK => clk, Q => n3682, QN
                           => n_1247);
   MY_CLK_r_REG1334_S1 : DFF_X1 port map( D => mult_143_n6204, CK => clk, Q => 
                           n3681, QN => n_1248);
   MY_CLK_r_REG1360_S1 : DFF_X1 port map( D => n1607, CK => clk, Q => n3680, QN
                           => n4614);
   MY_CLK_r_REG1361_S1 : DFF_X1 port map( D => mult_143_n1070, CK => clk, Q => 
                           n_1249, QN => n4615);
   MY_CLK_r_REG1259_S1 : DFF_X1 port map( D => n1604, CK => clk, Q => n3678, QN
                           => n4616);
   MY_CLK_r_REG1363_S1 : DFF_X1 port map( D => mult_143_n6174, CK => clk, Q => 
                           n3677, QN => n_1250);
   MY_CLK_r_REG1476_S1 : DFF_X1 port map( D => mult_143_n4407, CK => clk, Q => 
                           n3676, QN => n4617);
   MY_CLK_r_REG1493_S1 : DFF_X1 port map( D => mult_143_n2981, CK => clk, Q => 
                           n3675, QN => n4620);
   MY_CLK_r_REG1383_S1 : DFF_X1 port map( D => n1601, CK => clk, Q => n3674, QN
                           => n4619);
   MY_CLK_r_REG1423_S1 : DFF_X1 port map( D => mult_143_n4848, CK => clk, Q => 
                           n3673, QN => n_1251);
   MY_CLK_r_REG1410_S1 : DFF_X1 port map( D => mult_143_n5298, CK => clk, Q => 
                           n3672, QN => n4594);
   MY_CLK_r_REG1229_S2 : DFF_X1 port map( D => n1596, CK => clk, Q => n3670, QN
                           => n_1252);
   MY_CLK_r_REG1156_S2 : DFF_X1 port map( D => n3110, CK => clk, Q => n3669, QN
                           => n_1253);
   MY_CLK_r_REG1328_S2 : DFF_X1 port map( D => mult_143_n5258, CK => clk, Q => 
                           n3668, QN => n_1254);
   MY_CLK_r_REG1495_S1 : DFF_X1 port map( D => mult_143_n3443, CK => clk, Q => 
                           n3667, QN => n_1255);
   MY_CLK_r_REG1486_S1 : DFF_X1 port map( D => mult_143_n3137, CK => clk, Q => 
                           n3666, QN => n4595);
   MY_CLK_r_REG1498_S1 : DFF_X1 port map( D => mult_143_n3010, CK => clk, Q => 
                           n3665, QN => n4576);
   MY_CLK_r_REG1501_S1 : DFF_X1 port map( D => mult_143_n6626, CK => clk, Q => 
                           n3664, QN => n_1256);
   MY_CLK_r_REG1335_S1 : DFF_X1 port map( D => n1579, CK => clk, Q => n3663, QN
                           => n_1257);
   MY_CLK_r_REG1411_S1 : DFF_X1 port map( D => mult_143_n5310, CK => clk, Q => 
                           n3662, QN => n_1258);
   MY_CLK_r_REG1165_S2 : DFF_X1 port map( D => n1577, CK => clk, Q => n3660, QN
                           => n_1259);
   MY_CLK_r_REG1201_S1 : DFF_X1 port map( D => n1571, CK => clk, Q => n3658, QN
                           => n4577);
   MY_CLK_r_REG1505_S1 : DFF_X1 port map( D => n1061, CK => clk, Q => n3657, QN
                           => n_1260);
   MY_CLK_r_REG1504_S1 : DFF_X1 port map( D => mult_143_n3007, CK => clk, Q => 
                           n3656, QN => n_1261);
   MY_CLK_r_REG1491_S1 : DFF_X1 port map( D => mult_143_n6625, CK => clk, Q => 
                           n3655, QN => n_1262);
   MY_CLK_r_REG1473_S1 : DFF_X1 port map( D => n1071, CK => clk, Q => n3654, QN
                           => n_1263);
   MY_CLK_r_REG1488_S1 : DFF_X1 port map( D => n1565, CK => clk, Q => n3653, QN
                           => n_1264);
   MY_CLK_r_REG1489_S1 : DFF_X1 port map( D => n1075, CK => clk, Q => n3652, QN
                           => n_1265);
   MY_CLK_r_REG1370_S1 : DFF_X1 port map( D => n1564, CK => clk, Q => n3651, QN
                           => n_1266);
   MY_CLK_r_REG1484_S1 : DFF_X1 port map( D => n1085, CK => clk, Q => n3649, QN
                           => n4578);
   MY_CLK_r_REG1321_S1 : DFF_X1 port map( D => n571, CK => clk, Q => n3648, QN 
                           => n_1267);
   MY_CLK_r_REG1479_S1 : DFF_X1 port map( D => n1555, CK => clk, Q => n3647, QN
                           => n4597);
   MY_CLK_r_REG1316_S1 : DFF_X1 port map( D => mult_143_n74, CK => clk, Q => 
                           n3646, QN => n_1268);
   MY_CLK_r_REG1186_S3 : DFF_X1 port map( D => n2611, CK => clk, Q => n3642, QN
                           => n_1269);
   MY_CLK_r_REG1474_S1 : DFF_X1 port map( D => n1840, CK => clk, Q => n3641, QN
                           => n4596);
   MY_CLK_r_REG1462_S1 : DFF_X1 port map( D => n1756, CK => clk, Q => n3640, QN
                           => n_1270);
   MY_CLK_r_REG1461_S1 : DFF_X1 port map( D => n1754, CK => clk, Q => n3639, QN
                           => n_1271);
   MY_CLK_r_REG1440_S1 : DFF_X1 port map( D => n1741, CK => clk, Q => n3638, QN
                           => n_1272);
   MY_CLK_r_REG1442_S1 : DFF_X1 port map( D => n1742, CK => clk, Q => n3636, QN
                           => n_1273);
   MY_CLK_r_REG1420_S1 : DFF_X1 port map( D => n1719, CK => clk, Q => n3635, QN
                           => n_1274);
   MY_CLK_r_REG1418_S1 : DFF_X1 port map( D => n1745, CK => clk, Q => n3634, QN
                           => n_1275);
   MY_CLK_r_REG1315_S1 : DFF_X1 port map( D => n1730, CK => clk, Q => n3633, QN
                           => n_1276);
   MY_CLK_r_REG1312_S1 : DFF_X1 port map( D => n1736, CK => clk, Q => n3632, QN
                           => n_1277);
   MY_CLK_r_REG1313_S1 : DFF_X1 port map( D => n1734, CK => clk, Q => n3631, QN
                           => n_1278);
   MY_CLK_r_REG1314_S1 : DFF_X1 port map( D => n1733, CK => clk, Q => n3630, QN
                           => n_1279);
   MY_CLK_r_REG1149_S1 : DFF_X1 port map( D => n1727, CK => clk, Q => n3629, QN
                           => n_1280);
   MY_CLK_r_REG1197_S1 : DFF_X1 port map( D => n1737, CK => clk, Q => n3628, QN
                           => n_1281);
   MY_CLK_r_REG1168_S1 : DFF_X1 port map( D => n1735, CK => clk, Q => n3627, QN
                           => n_1282);
   MY_CLK_r_REG1342_S1 : DFF_X1 port map( D => n1729, CK => clk, Q => n3626, QN
                           => n_1283);
   MY_CLK_r_REG1392_S1 : DFF_X1 port map( D => n2709, CK => clk, Q => n3625, QN
                           => n_1284);
   MY_CLK_r_REG1414_S1 : DFF_X1 port map( D => n1748, CK => clk, Q => n3624, QN
                           => n_1285);
   MY_CLK_r_REG1408_S1 : DFF_X1 port map( D => n1720, CK => clk, Q => n3623, QN
                           => n_1286);
   MY_CLK_r_REG1409_S1 : DFF_X1 port map( D => n2746, CK => clk, Q => n3622, QN
                           => n_1287);
   MY_CLK_r_REG1390_S1 : DFF_X1 port map( D => n1744, CK => clk, Q => n3621, QN
                           => n_1288);
   MY_CLK_r_REG1384_S1 : DFF_X1 port map( D => n1751, CK => clk, Q => n3620, QN
                           => n_1289);
   MY_CLK_r_REG1341_S1 : DFF_X1 port map( D => n1732, CK => clk, Q => n3619, QN
                           => n_1290);
   MY_CLK_r_REG1435_S1 : DFF_X1 port map( D => n1721, CK => clk, Q => n3618, QN
                           => n_1291);
   MY_CLK_r_REG1436_S1 : DFF_X1 port map( D => n1753, CK => clk, Q => n3617, QN
                           => n_1292);
   MY_CLK_r_REG1437_S1 : DFF_X1 port map( D => n1743, CK => clk, Q => n3616, QN
                           => n_1293);
   MY_CLK_r_REG1438_S1 : DFF_X1 port map( D => n1746, CK => clk, Q => n3615, QN
                           => n_1294);
   MY_CLK_r_REG1212_S3 : DFF_X1 port map( D => n1750, CK => clk, Q => n3614, QN
                           => n_1295);
   MY_CLK_r_REG1481_S1 : DFF_X1 port map( D => n1582, CK => clk, Q => n3613, QN
                           => n_1296);
   MY_CLK_r_REG1227_S2 : DFF_X1 port map( D => mult_143_n5468, CK => clk, Q => 
                           n3610, QN => n4854);
   MY_CLK_r_REG1308_S2 : DFF_X1 port map( D => n1634, CK => clk, Q => n3609, QN
                           => n_1297);
   MY_CLK_r_REG1153_S2 : DFF_X1 port map( D => mult_143_n5397, CK => clk, Q => 
                           n3608, QN => n4722);
   MY_CLK_r_REG1299_S2 : DFF_X1 port map( D => n2972, CK => clk, Q => n_1298, 
                           QN => n4906);
   MY_CLK_r_REG1162_S2 : DFF_X1 port map( D => n1680, CK => clk, Q => n3605, QN
                           => n_1299);
   MY_CLK_r_REG1237_S2 : DFF_X1 port map( D => n2987, CK => clk, Q => n3603, QN
                           => n_1300);
   MY_CLK_r_REG1306_S2 : DFF_X1 port map( D => n1570, CK => clk, Q => n3602, QN
                           => n_1301);
   MY_CLK_r_REG1330_S2 : DFF_X1 port map( D => mult_143_n5257, CK => clk, Q => 
                           n3601, QN => n_1302);
   MY_CLK_r_REG1171_S2 : DFF_X1 port map( D => n3026, CK => clk, Q => n3598, QN
                           => n4862);
   MY_CLK_r_REG1451_S1 : DFF_X1 port map( D => mult_143_n5859, CK => clk, Q => 
                           n3597, QN => n4591);
   MY_CLK_r_REG1353_S1 : DFF_X1 port map( D => mult_143_n4824, CK => clk, Q => 
                           n3596, QN => n_1303);
   MY_CLK_r_REG1300_S2 : DFF_X1 port map( D => mult_143_n5394, CK => clk, Q => 
                           n3595, QN => n_1304);
   MY_CLK_r_REG1141_S2 : DFF_X1 port map( D => n4864, CK => clk, Q => n3593, QN
                           => n_1305);
   MY_CLK_r_REG1157_S2 : DFF_X1 port map( D => n3110, CK => clk, Q => n3592, QN
                           => n_1306);
   MY_CLK_r_REG1217_S2 : DFF_X1 port map( D => n1638, CK => clk, Q => n3591, QN
                           => n_1307);
   MY_CLK_r_REG1258_S1 : DFF_X1 port map( D => n993, CK => clk, Q => n3590, QN 
                           => n4593);
   MY_CLK_r_REG1256_S1 : DFF_X1 port map( D => n1549, CK => clk, Q => n3589, QN
                           => n4579);
   MY_CLK_r_REG1255_S1 : DFF_X1 port map( D => n1548, CK => clk, Q => n3588, QN
                           => n4580);
   MY_CLK_r_REG1460_S1 : DFF_X1 port map( D => mult_143_n5817, CK => clk, Q => 
                           n3587, QN => n_1308);
   MY_CLK_r_REG1447_S1 : DFF_X1 port map( D => mult_143_n5884, CK => clk, Q => 
                           n3586, QN => n_1309);
   MY_CLK_r_REG1459_S1 : DFF_X1 port map( D => mult_143_n5823, CK => clk, Q => 
                           n3585, QN => n_1310);
   MY_CLK_r_REG1458_S1 : DFF_X1 port map( D => mult_143_n5808, CK => clk, Q => 
                           n3584, QN => n_1311);
   MY_CLK_r_REG1448_S1 : DFF_X1 port map( D => mult_143_n5875, CK => clk, Q => 
                           n3583, QN => n_1312);
   MY_CLK_r_REG1422_S1 : DFF_X1 port map( D => mult_143_n5926, CK => clk, Q => 
                           n3582, QN => n_1313);
   MY_CLK_r_REG1396_S1 : DFF_X1 port map( D => mult_143_n5963, CK => clk, Q => 
                           n3581, QN => n_1314);
   MY_CLK_r_REG1169_S1 : DFF_X1 port map( D => mult_143_n6074, CK => clk, Q => 
                           n3580, QN => n_1315);
   MY_CLK_r_REG1455_S1 : DFF_X1 port map( D => n1544, CK => clk, Q => n3579, QN
                           => n_1316);
   MY_CLK_r_REG1421_S1 : DFF_X1 port map( D => mult_143_n5929, CK => clk, Q => 
                           n3578, QN => n_1317);
   MY_CLK_r_REG1124_S3 : DFF_X1 port map( D => mult_143_n4776, CK => clk, Q => 
                           n3577, QN => n_1318);
   MY_CLK_r_REG1347_S1 : DFF_X1 port map( D => mult_143_n6037, CK => clk, Q => 
                           n3576, QN => n_1319);
   MY_CLK_r_REG1346_S1 : DFF_X1 port map( D => mult_143_n6015, CK => clk, Q => 
                           n3575, QN => n_1320);
   MY_CLK_r_REG1456_S1 : DFF_X1 port map( D => mult_143_n5820, CK => clk, Q => 
                           n3574, QN => n_1321);
   MY_CLK_r_REG1449_S1 : DFF_X1 port map( D => mult_143_n5881, CK => clk, Q => 
                           n3573, QN => n_1322);
   MY_CLK_r_REG1445_S1 : DFF_X1 port map( D => mult_143_n6195, CK => clk, Q => 
                           n3572, QN => n_1323);
   MY_CLK_r_REG1344_S1 : DFF_X1 port map( D => mult_143_n6018, CK => clk, Q => 
                           n3571, QN => n_1324);
   MY_CLK_r_REG1345_S1 : DFF_X1 port map( D => mult_143_n4893, CK => clk, Q => 
                           n3570, QN => n_1325);
   MY_CLK_r_REG1417_S1 : DFF_X1 port map( D => mult_143_n6250, CK => clk, Q => 
                           n3569, QN => n_1326);
   MY_CLK_r_REG1394_S1 : DFF_X1 port map( D => mult_143_n4826, CK => clk, Q => 
                           n3568, QN => n_1327);
   MY_CLK_r_REG1250_S1 : DFF_X1 port map( D => n1535, CK => clk, Q => n3567, QN
                           => n4604);
   MY_CLK_r_REG1254_S1 : DFF_X1 port map( D => n1534, CK => clk, Q => n3566, QN
                           => n4605);
   MY_CLK_r_REG1318_S1 : DFF_X1 port map( D => mult_143_n4934, CK => clk, Q => 
                           n3565, QN => n_1328);
   MY_CLK_r_REG1249_S1 : DFF_X1 port map( D => n1533, CK => clk, Q => n3564, QN
                           => n4606);
   MY_CLK_r_REG1187_S1 : DFF_X1 port map( D => mult_143_n4931, CK => clk, Q => 
                           n3563, QN => n_1329);
   MY_CLK_r_REG1446_S1 : DFF_X1 port map( D => mult_143_n5900, CK => clk, Q => 
                           n3562, QN => n_1330);
   MY_CLK_r_REG1399_S1 : DFF_X1 port map( D => mult_143_n5981, CK => clk, Q => 
                           n3561, QN => n_1331);
   MY_CLK_r_REG1419_S1 : DFF_X1 port map( D => n1524, CK => clk, Q => n3560, QN
                           => n_1332);
   MY_CLK_r_REG1302_S1 : DFF_X1 port map( D => n1522, CK => clk, Q => n3559, QN
                           => n_1333);
   MY_CLK_r_REG1377_S1 : DFF_X1 port map( D => mult_143_n6169, CK => clk, Q => 
                           n3558, QN => n_1334);
   MY_CLK_r_REG1403_S1 : DFF_X1 port map( D => mult_143_n1101, CK => clk, Q => 
                           n_1335, QN => n4608);
   MY_CLK_r_REG1323_S1 : DFF_X1 port map( D => mult_143_n4962, CK => clk, Q => 
                           n3556, QN => n_1336);
   MY_CLK_r_REG1234_S2 : DFF_X1 port map( D => n1517, CK => clk, Q => n3555, QN
                           => n4609);
   MY_CLK_r_REG1369_S1 : DFF_X1 port map( D => mult_143_n5192, CK => clk, Q => 
                           n3552, QN => n_1337);
   MY_CLK_r_REG1175_S1 : DFF_X1 port map( D => n1515, CK => clk, Q => n3551, QN
                           => n_1338);
   MY_CLK_r_REG1317_S1 : DFF_X1 port map( D => mult_143_n4886, CK => clk, Q => 
                           n_1339, QN => n4751);
   MY_CLK_r_REG1395_S1 : DFF_X1 port map( D => mult_143_n6239, CK => clk, Q => 
                           n4894, QN => n_1340);
   MY_CLK_r_REG1144_S2 : DFF_X1 port map( D => n1508, CK => clk, Q => n3548, QN
                           => n4879);
   MY_CLK_r_REG1322_S1 : DFF_X1 port map( D => mult_143_n5195, CK => clk, Q => 
                           n3547, QN => n_1341);
   MY_CLK_r_REG1349_S1 : DFF_X1 port map( D => n1505, CK => clk, Q => n3546, QN
                           => n_1342);
   MY_CLK_r_REG1348_S1 : DFF_X1 port map( D => mult_143_n4876, CK => clk, Q => 
                           n3545, QN => n_1343);
   MY_CLK_r_REG1042_S3 : DFF_X1 port map( D => n385, CK => clk, Q => n3544, QN 
                           => n_1344);
   MY_CLK_r_REG1350_S1 : DFF_X1 port map( D => n1500, CK => clk, Q => n3543, QN
                           => n_1345);
   MY_CLK_r_REG1374_S1 : DFF_X1 port map( D => mult_143_n4942, CK => clk, Q => 
                           n3542, QN => n_1346);
   MY_CLK_r_REG1351_S1 : DFF_X1 port map( D => n1499, CK => clk, Q => n3541, QN
                           => n_1347);
   MY_CLK_r_REG1397_S1 : DFF_X1 port map( D => mult_143_n48, CK => clk, Q => 
                           n3538, QN => n_1348);
   MY_CLK_r_REG1424_S1 : DFF_X1 port map( D => mult_143_n36, CK => clk, Q => 
                           n3537, QN => n_1349);
   MY_CLK_r_REG1126_S3 : DFF_X1 port map( D => mult_143_n4771, CK => clk, Q => 
                           n3535, QN => n_1350);
   MY_CLK_r_REG1354_S1 : DFF_X1 port map( D => mult_143_n72, CK => clk, Q => 
                           n3533, QN => n_1351);
   MY_CLK_r_REG1464_S1 : DFF_X1 port map( D => mult_143_n5811, CK => clk, Q => 
                           n3532, QN => n_1352);
   MY_CLK_r_REG1467_S1 : DFF_X1 port map( D => mult_143_n5831, CK => clk, Q => 
                           n3530, QN => n_1353);
   MY_CLK_r_REG1398_S1 : DFF_X1 port map( D => mult_143_n5979, CK => clk, Q => 
                           n3529, QN => n_1354);
   MY_CLK_r_REG1352_S1 : DFF_X1 port map( D => mult_143_n6034, CK => clk, Q => 
                           n3528, QN => n_1355);
   MY_CLK_r_REG1039_S1 : DFF_X1 port map( D => mult_143_n4851, CK => clk, Q => 
                           n3526, QN => n_1356);
   MY_CLK_r_REG1320_S1 : DFF_X1 port map( D => mult_143_n4988, CK => clk, Q => 
                           n3525, QN => n_1357);
   MY_CLK_r_REG1180_S2 : DFF_X1 port map( D => n1476, CK => clk, Q => n3524, QN
                           => n_1358);
   MY_CLK_r_REG1179_S2 : DFF_X1 port map( D => mult_143_n5699, CK => clk, Q => 
                           n3523, QN => n_1359);
   MY_CLK_r_REG1362_S1 : DFF_X1 port map( D => mult_143_n6282, CK => clk, Q => 
                           n_1360, QN => n4956);
   MY_CLK_r_REG1158_S1 : DFF_X1 port map( D => mult_143_n4913, CK => clk, Q => 
                           n3521, QN => n_1361);
   MY_CLK_r_REG1304_S1 : DFF_X1 port map( D => mult_143_n6261, CK => clk, Q => 
                           n3520, QN => n_1362);
   MY_CLK_r_REG1432_S1 : DFF_X1 port map( D => mult_143_n5119, CK => clk, Q => 
                           n3519, QN => n_1363);
   MY_CLK_r_REG1472_S1 : DFF_X1 port map( D => mult_143_n6120, CK => clk, Q => 
                           n3518, QN => n4771);
   MY_CLK_r_REG1444_S1 : DFF_X1 port map( D => mult_143_n2334, CK => clk, Q => 
                           n3517, QN => n_1364);
   MY_CLK_r_REG1508_S1 : DFF_X1 port map( D => mult_143_n1818, CK => clk, Q => 
                           n3516, QN => n_1365);
   MY_CLK_r_REG1239_S2 : DFF_X1 port map( D => n1494, CK => clk, Q => n3515, QN
                           => n_1366);
   MY_CLK_r_REG1310_S2 : DFF_X1 port map( D => mult_143_n5372, CK => clk, Q => 
                           n_1367, QN => n4905);
   MY_CLK_r_REG1160_S2 : DFF_X1 port map( D => n1493, CK => clk, Q => n3513, QN
                           => n_1368);
   MY_CLK_r_REG1222_S2 : DFF_X1 port map( D => n1491, CK => clk, Q => n3512, QN
                           => n_1369);
   MY_CLK_r_REG1216_S2 : DFF_X1 port map( D => n1490, CK => clk, Q => n3511, QN
                           => n_1370);
   MY_CLK_r_REG1150_S2 : DFF_X1 port map( D => n1489, CK => clk, Q => n3510, QN
                           => n_1371);
   MY_CLK_r_REG1307_S2 : DFF_X1 port map( D => n1484, CK => clk, Q => n3508, QN
                           => n4573);
   MY_CLK_r_REG1305_S2 : DFF_X1 port map( D => n1483, CK => clk, Q => n3507, QN
                           => n_1372);
   MY_CLK_r_REG1203_S2 : DFF_X1 port map( D => mult_143_n5424, CK => clk, Q => 
                           n3505, QN => n_1373);
   MY_CLK_r_REG1260_S1 : DFF_X1 port map( D => n1481, CK => clk, Q => n3504, QN
                           => n_1374);
   MY_CLK_r_REG1331_S2 : DFF_X1 port map( D => n1479, CK => clk, Q => n3502, QN
                           => n_1375);
   MY_CLK_r_REG1226_S2 : DFF_X1 port map( D => mult_143_n5469, CK => clk, Q => 
                           n3499, QN => n_1376);
   MY_CLK_r_REG1155_S2 : DFF_X1 port map( D => n1067, CK => clk, Q => n3496, QN
                           => n4896);
   MY_CLK_r_REG1173_S2 : DFF_X1 port map( D => n2924, CK => clk, Q => n3495, QN
                           => n_1377);
   MY_CLK_r_REG1161_S2 : DFF_X1 port map( D => n1470, CK => clk, Q => n3494, QN
                           => n4829);
   MY_CLK_r_REG1174_S2 : DFF_X1 port map( D => n2924, CK => clk, Q => n3492, QN
                           => n4716);
   MY_CLK_r_REG1233_S2 : DFF_X1 port map( D => mult_143_n5730, CK => clk, Q => 
                           n3490, QN => n_1378);
   MY_CLK_r_REG1142_S2 : DFF_X1 port map( D => mult_143_n5574, CK => clk, Q => 
                           n3489, QN => n4904);
   U1500 : INV_X1 port map( A => n1647, ZN => n2672);
   U1501 : INV_X1 port map( A => n1689, ZN => n2767);
   U1502 : INV_X1 port map( A => n1573, ZN => n2686);
   U1504 : INV_X1 port map( A => n1568, ZN => n2688);
   U1505 : INV_X1 port map( A => n1712, ZN => n2762);
   U1507 : INV_X1 port map( A => n3120, ZN => n2605);
   U1509 : INV_X1 port map( A => n1673, ZN => n2718);
   U1512 : INV_X1 port map( A => n1556, ZN => n2690);
   U1517 : INV_X1 port map( A => n1631, ZN => n2782);
   U1523 : INV_X1 port map( A => n1574, ZN => n2685);
   U1526 : INV_X1 port map( A => n4760, ZN => n2749);
   U1527 : INV_X1 port map( A => n1488, ZN => n2713);
   U1540 : INV_X1 port map( A => n1731, ZN => n2689);
   U1546 : INV_X1 port map( A => n1651, ZN => n2703);
   U1556 : INV_X1 port map( A => B_SIG(12), ZN => n2841);
   U1564 : INV_X1 port map( A => mult_143_n4959, ZN => n2706);
   U1577 : INV_X1 port map( A => mult_143_n5899, ZN => n2811);
   n1724 <= '1';
   U1503 : INV_X1 port map( A => n1657, ZN => n2695);
   U1445 : AOI222_X1 port map( A1 => n4886, A2 => mult_143_n5556, B1 => 
                           mult_143_n5556, B2 => mult_143_n5554, C1 => 
                           mult_143_n5557, C2 => mult_143_n5554, ZN => 
                           mult_143_n5395);
   MY_CLK_r_REG1490_S1 : DFF_X2 port map( D => B_SIG(16), CK => clk, Q => n3783
                           , QN => n4746);
   MY_CLK_r_REG1471_S1 : DFF_X1 port map( D => B_SIG(23), CK => clk, Q => n3790
                           , QN => n4770);
   MY_CLK_r_REG1492_S1 : DFF_X1 port map( D => B_SIG(15), CK => clk, Q => n3782
                           , QN => n4761);
   MY_CLK_r_REG1332_S1 : DFF_X1 port map( D => A_SIG(17), CK => clk, Q => n3796
                           , QN => n4759);
   MY_CLK_r_REG1391_S1 : DFF_X1 port map( D => n1765, CK => clk, Q => n3774, QN
                           => n4753);
   MY_CLK_r_REG1303_S1 : DFF_X1 port map( D => A_SIG(20), CK => clk, Q => n3797
                           , QN => n4749);
   MY_CLK_r_REG1485_S1 : DFF_X1 port map( D => B_SIG(18), CK => clk, Q => n3785
                           , QN => n4748);
   MY_CLK_r_REG1480_S1 : DFF_X2 port map( D => B_SIG(20), CK => clk, Q => n3787
                           , QN => n4681);
   MY_CLK_r_REG1325_S1 : DFF_X1 port map( D => mult_143_n4842, CK => clk, Q => 
                           n3645, QN => n4672);
   MY_CLK_r_REG1439_S1 : DFF_X1 port map( D => n642, CK => clk, Q => n3768, QN 
                           => n4721);
   MY_CLK_r_REG1154_S2 : DFF_X1 port map( D => n3010, CK => clk, Q => n3600, QN
                           => n_1379);
   MY_CLK_r_REG1151_S2 : DFF_X1 port map( D => mult_143_n5393, CK => clk, Q => 
                           n3606, QN => n_1380);
   MY_CLK_r_REG1468_S1 : DFF_X1 port map( D => n536, CK => clk, Q => n3769, QN 
                           => n4730);
   MY_CLK_r_REG1176_S2 : DFF_X1 port map( D => mult_143_n5680, CK => clk, Q => 
                           n3671, QN => n_1381);
   MY_CLK_r_REG1494_S1 : DFF_X1 port map( D => B_SIG(14), CK => clk, Q => n3781
                           , QN => n4735);
   MY_CLK_r_REG1248_S1 : DFF_X1 port map( D => n748, CK => clk, Q => n3775, QN 
                           => n4752);
   MY_CLK_r_REG1380_S1 : DFF_X1 port map( D => A_SIG(11), CK => clk, Q => n3794
                           , QN => n4768);
   MY_CLK_r_REG1167_S1 : DFF_X1 port map( D => n2598, CK => clk, Q => n3772, QN
                           => n4676);
   mult_143_U3441 : NOR2_X2 port map( A1 => A_SIG(0), A2 => n639, ZN => 
                           mult_143_n3245);
   U360 : NAND2_X1 port map( A1 => n629, A2 => B_SIG(1), ZN => mult_143_n6302);
   U206 : INV_X2 port map( A => n4752, ZN => n2840);
   U838 : OR2_X1 port map( A1 => n4599, A2 => n4604, ZN => n2691);
   mult_143_U3784 : NAND2_X1 port map( A1 => n3790, A2 => n3518, ZN => n1589);
   U169 : XNOR2_X1 port map( A => n910, B => mult_143_n6302, ZN => n2817);
   mult_143_U3443 : NOR2_X2 port map( A1 => mult_143_n5853, A2 => n638, ZN => 
                           mult_143_n2);
   mult_143_U3054 : NOR2_X1 port map( A1 => mult_143_n5484, A2 => 
                           mult_143_n5485, ZN => n984);
   U1259 : INV_X1 port map( A => n979, ZN => n804);
   U275 : AOI21_X1 port map( B1 => n812, B2 => mult_143_n6078, A => 
                           mult_143_n6080, ZN => mult_143_n5970);
   U1193 : AOI222_X1 port map( A1 => n3818, A2 => n1647, B1 => n3818, B2 => 
                           n3707, C1 => n1647, C2 => n3707, ZN => 
                           mult_143_n5439);
   U4 : OR2_X1 port map( A1 => mult_143_n5153, A2 => mult_143_n5152, ZN => 
                           mult_143_n4401);
   MY_CLK_r_REG1329_S2 : DFF_X1 port map( D => mult_143_n5255, CK => clk, Q => 
                           n3554, QN => n_1382);
   MY_CLK_r_REG1301_S2 : DFF_X1 port map( D => mult_143_n5395, CK => clk, Q => 
                           n3488, QN => n_1383);
   MY_CLK_r_REG1219_S2 : DFF_X1 port map( D => n4729, CK => clk, Q => n3501, QN
                           => n_1384);
   MY_CLK_r_REG1228_S2 : DFF_X1 port map( D => n2980, CK => clk, Q => n_1385, 
                           QN => n4963);
   MY_CLK_r_REG1404_S1 : DFF_X1 port map( D => n1747, CK => clk, Q => n3612, QN
                           => n_1386);
   MY_CLK_r_REG1190_S2 : DFF_X1 port map( D => n1486, CK => clk, Q => n3509, QN
                           => n4570);
   MY_CLK_r_REG1385_S1 : DFF_X1 port map( D => mult_143_n5320, CK => clk, Q => 
                           n3726, QN => n_1387);
   MY_CLK_r_REG1244_S2 : DFF_X1 port map( D => n1714, CK => clk, Q => n3760, QN
                           => n_1388);
   MY_CLK_r_REG1117_S3 : DFF_X1 port map( D => n2947, CK => clk, Q => n3776, QN
                           => n_1389);
   U5 : INV_X1 port map( A => n4735, ZN => n4736);
   U15 : AOI222_X1 port map( A1 => n3610, A2 => n3829, B1 => n3610, B2 => n3499
                           , C1 => n3829, C2 => n3499, ZN => n1474);
   U28 : XNOR2_X1 port map( A => mult_143_n809, B => n4713, ZN => 
                           mult_143_n5647);
   U35 : NAND2_X1 port map( A1 => n4647, A2 => n4628, ZN => mult_143_n5707);
   U46 : XNOR2_X1 port map( A => n2627, B => n4788, ZN => mult_143_n5760);
   U60 : XNOR2_X1 port map( A => n4821, B => n3064, ZN => mult_143_n5708);
   U69 : XNOR2_X1 port map( A => n2732, B => n4795, ZN => mult_143_n5531);
   U100 : OR2_X1 port map( A1 => n4775, A2 => n4774, ZN => mult_143_n5163);
   U111 : XNOR2_X1 port map( A => mult_143_n5611, B => n4607, ZN => 
                           mult_143_n5419);
   U113 : XNOR2_X1 port map( A => mult_143_n5896, B => n3099, ZN => n2730);
   U127 : NOR2_X1 port map( A1 => mult_143_n5090, A2 => n436, ZN => 
                           mult_143_n5089);
   U134 : NOR2_X1 port map( A1 => n4645, A2 => n569, ZN => n568);
   U143 : OR2_X1 port map( A1 => n403, A2 => n4808, ZN => n4807);
   U168 : XNOR2_X1 port map( A => n1474, B => n4640, ZN => mult_143_n5437);
   U194 : XNOR2_X1 port map( A => n3599, B => n3708, ZN => n1645);
   U227 : AND2_X1 port map( A1 => n3784, A2 => n3819, ZN => n4644);
   U232 : XNOR2_X1 port map( A => n3751, B => n3524, ZN => n4641);
   U255 : NOR2_X1 port map( A1 => n3643, A2 => n4596, ZN => n4808);
   U289 : NOR2_X1 port map( A1 => mult_143_n5443, A2 => n4644, ZN => n1516);
   U293 : CLKBUF_X1 port map( A => mult_143_n4768, Z => n3117);
   U298 : AOI222_X1 port map( A1 => n4762, A2 => n3733, B1 => n4762, B2 => 
                           n3734, C1 => n3733, C2 => n3734, ZN => 
                           mult_143_n5207);
   U343 : INV_X1 port map( A => mult_143_n1017, ZN => n2711);
   U367 : INV_X1 port map( A => n4681, ZN => n2908);
   U379 : AOI222_X1 port map( A1 => n2632, A2 => n4588, B1 => n4843, B2 => 
                           n2632, C1 => n2799, C2 => n4588, ZN => 
                           mult_143_n5346);
   U405 : XNOR2_X1 port map( A => n1597, B => n3696, ZN => n4640);
   U475 : OR2_X1 port map( A1 => n4601, A2 => mult_143_n1898, ZN => n2667);
   U477 : XNOR2_X1 port map( A => n2667, B => n4789, ZN => n4788);
   U486 : OAI221_X1 port map( B1 => n3511, B2 => n4637, C1 => n4639, C2 => 
                           mult_143_n5516, A => mult_143_n5221, ZN => n944);
   U507 : AOI222_X1 port map( A1 => n2812, A2 => n3112, B1 => n2812, B2 => 
                           n2679, C1 => n3112, C2 => n2679, ZN => 
                           mult_143_n5477);
   U523 : XOR2_X1 port map( A => n4602, B => mult_143_n5610, Z => 
                           mult_143_n5420);
   U527 : INV_X2 port map( A => n4632, ZN => mult_143_n4490);
   U528 : OR2_X1 port map( A1 => n4634, A2 => n2780, ZN => n2631);
   U646 : AOI222_X1 port map( A1 => mult_143_n5559, A2 => n2756, B1 => 
                           mult_143_n5561, B2 => mult_143_n5559, C1 => n2756, 
                           C2 => mult_143_n5561, ZN => mult_143_n5401);
   U691 : OAI22_X1 port map( A1 => mult_143_n5163, A2 => n4790, B1 => 
                           mult_143_n5164, B2 => n3106, ZN => mult_143_n5184);
   U700 : NOR2_X1 port map( A1 => mult_143_n6097, A2 => mult_143_n6098, ZN => 
                           mult_143_n6040);
   U717 : XNOR2_X1 port map( A => mult_143_n5647, B => n4642, ZN => n1051);
   U734 : XNOR2_X1 port map( A => n4809, B => n975, ZN => mult_143_n5796);
   U747 : CLKBUF_X1 port map( A => A_SIG(23), Z => n748);
   U753 : NAND2_X1 port map( A1 => n651, A2 => mult_143_n6300, ZN => 
                           mult_143_n4842);
   U758 : CLKBUF_X1 port map( A => mult_143_n76, Z => n1027);
   U772 : OR2_X1 port map( A1 => mult_143_n5440, A2 => mult_143_n5441, ZN => 
                           n4567);
   U783 : OR2_X1 port map( A1 => n1624, A2 => n1625, ZN => n4569);
   U787 : OR2_X1 port map( A1 => mult_143_n5505, A2 => mult_143_n5508, ZN => 
                           n4574);
   U790 : XNOR2_X1 port map( A => n3803, B => n3582, ZN => n4583);
   U796 : XOR2_X1 port map( A => n3775, B => n3580, Z => n4585);
   U799 : XOR2_X1 port map( A => n3576, B => n4760, Z => n4586);
   U801 : XNOR2_X1 port map( A => n3769, B => n3574, ZN => n4587);
   U802 : XNOR2_X1 port map( A => n3768, B => n3573, ZN => n4588);
   U804 : OR2_X1 port map( A1 => n3645, A2 => n3655, ZN => n4598);
   U814 : OR2_X1 port map( A1 => mult_143_n5288, A2 => mult_143_n5289, ZN => 
                           n4600);
   U828 : XOR2_X1 port map( A => n4760, B => n3571, Z => n4602);
   U834 : XNOR2_X1 port map( A => n3774, B => n1503, ZN => n4607);
   U848 : XNOR2_X1 port map( A => n3769, B => n3532, ZN => n4611);
   U857 : XNOR2_X1 port map( A => mult_143_n6148, B => mult_143_n6149, ZN => 
                           n4623);
   U867 : OR2_X1 port map( A1 => n2719, A2 => mult_143_n6367, ZN => n4628);
   U881 : INV_X1 port map( A => mult_143_n1898, ZN => n1551);
   U905 : INV_X1 port map( A => mult_143_n1902, ZN => n1550);
   U914 : INV_X1 port map( A => mult_143_n1900, ZN => n1552);
   U916 : XNOR2_X1 port map( A => n3695, B => n3526, ZN => n4633);
   U926 : OR2_X1 port map( A1 => n2726, A2 => n3795, ZN => n4635);
   U963 : XOR2_X1 port map( A => n2840, B => mult_143_n6086, Z => n4638);
   U967 : INV_X1 port map( A => mult_143_n5648, ZN => n4642);
   U972 : INV_X1 port map( A => n4769, ZN => n1584);
   U991 : XNOR2_X1 port map( A => n1645, B => n4641, ZN => mult_143_n5696);
   U993 : NAND2_X1 port map( A1 => n4598, A2 => n4646, ZN => n4645);
   U1000 : INV_X1 port map( A => n4737, ZN => n4646);
   U1012 : INV_X1 port map( A => mult_143_n777, ZN => mult_143_n6563);
   U1014 : NAND2_X1 port map( A1 => mult_143_n777, A2 => n4648, ZN => n4647);
   U1018 : NAND2_X1 port map( A1 => n2719, A2 => mult_143_n6367, ZN => n4648);
   U1020 : NOR2_X1 port map( A1 => n4649, A2 => n3034, ZN => n4819);
   U1025 : XOR2_X1 port map( A => n3118, B => n2835, Z => n4649);
   U1026 : XOR2_X1 port map( A => mult_143_n4994, B => mult_143_n4995, Z => 
                           n4650);
   U1027 : OR2_X1 port map( A1 => n2982, A2 => n2981, ZN => mult_143_n5683);
   U1035 : XNOR2_X1 port map( A => mult_143_n5089, B => n4752, ZN => n4651);
   U1040 : XOR2_X1 port map( A => mult_143_n5087, B => mult_143_n5086, Z => 
                           n4652);
   U1041 : XOR2_X1 port map( A => mult_143_n5087, B => mult_143_n5086, Z => 
                           n3048);
   U1042 : AOI222_X1 port map( A1 => n2715, A2 => mult_143_n5462, B1 => n2715, 
                           B2 => mult_143_n5463, C1 => mult_143_n5462, C2 => 
                           mult_143_n5463, ZN => n4653);
   U1061 : OAI21_X1 port map( B1 => mult_143_n5435, B2 => mult_143_n5434, A => 
                           mult_143_n3075, ZN => mult_143_n5432);
   U1066 : XNOR2_X1 port map( A => n4638, B => n2895, ZN => n4798);
   U1075 : INV_X1 port map( A => n4692, ZN => n4656);
   U1084 : XOR2_X1 port map( A => n4657, B => n3578, Z => n1731);
   U1085 : XNOR2_X1 port map( A => mult_143_n4944, B => n3774, ZN => n4658);
   U1089 : XNOR2_X1 port map( A => mult_143_n4944, B => n3774, ZN => 
                           mult_143_n4939);
   U1105 : XNOR2_X1 port map( A => mult_143_n4915, B => n4661, ZN => n2610);
   U1117 : XNOR2_X1 port map( A => n1625, B => n1624, ZN => n4661);
   U1130 : AOI222_X1 port map( A1 => n2610, A2 => n4671, B1 => n2610, B2 => 
                           mult_143_n5178, C1 => mult_143_n5177, C2 => 
                           mult_143_n5178, ZN => n4662);
   U1143 : AOI222_X1 port map( A1 => n2610, A2 => n4671, B1 => n2610, B2 => 
                           mult_143_n5178, C1 => mult_143_n5177, C2 => 
                           mult_143_n5178, ZN => mult_143_n5160);
   U1145 : AND2_X1 port map( A1 => mult_143_n5181, A2 => mult_143_n5182, ZN => 
                           n4801);
   U1153 : XNOR2_X1 port map( A => n3759, B => n3683, ZN => mult_143_n5309);
   U1159 : INV_X1 port map( A => n4719, ZN => n4664);
   U1182 : AOI222_X1 port map( A1 => mult_143_n5067, A2 => n3803, B1 => 
                           mult_143_n5067, B2 => n667, C1 => n3803, C2 => n667,
                           ZN => mult_143_n686);
   U1195 : AOI222_X1 port map( A1 => mult_143_n4939, A2 => n4630, B1 => 
                           mult_143_n4939, B2 => mult_143_n4937, C1 => 
                           mult_143_n4937, C2 => n4630, ZN => n4669);
   U1208 : INV_X1 port map( A => n4730, ZN => n4670);
   U1209 : XNOR2_X1 port map( A => mult_143_n5416, B => n2691, ZN => n4671);
   U1211 : XOR2_X1 port map( A => mult_143_n917, B => n3062, Z => 
                           mult_143_n5623);
   U1214 : NAND2_X1 port map( A1 => n3024, A2 => n2636, ZN => n4673);
   U1216 : OAI21_X1 port map( B1 => n3130, B2 => mult_143_n4915, A => n4569, ZN
                           => n965);
   U1220 : XNOR2_X1 port map( A => n3118, B => n2835, ZN => n4674);
   U1224 : INV_X1 port map( A => n4761, ZN => n4675);
   U1229 : INV_X1 port map( A => n4676, ZN => n4677);
   U1236 : OAI22_X1 port map( A1 => n4679, A2 => n4629, B1 => n4680, B2 => 
                           n4770, ZN => n4678);
   U1250 : XNOR2_X1 port map( A => n1670, B => n4780, ZN => n2766);
   U1252 : XNOR2_X1 port map( A => mult_143_n5765, B => n4682, ZN => 
                           mult_143_n5466);
   U1261 : XOR2_X1 port map( A => mult_143_n686, B => mult_143_n6348, Z => 
                           n4682);
   U1274 : XNOR2_X1 port map( A => mult_143_n5566, B => mult_143_n5604, ZN => 
                           mult_143_n5561);
   U1279 : XNOR2_X1 port map( A => n2704, B => n4683, ZN => mult_143_n5701);
   U1281 : XNOR2_X1 port map( A => mult_143_n6361, B => mult_143_n6362, ZN => 
                           n4683);
   U1349 : XNOR2_X1 port map( A => mult_143_n5387, B => n2888, ZN => n4686);
   U1366 : AOI222_X1 port map( A1 => mult_143_n6427, A2 => n2877, B1 => 
                           mult_143_n6427, B2 => n2705, C1 => n2877, C2 => 
                           n2705, ZN => mult_143_n5389);
   U1375 : AOI222_X1 port map( A1 => n3047, A2 => mult_143_n5625, B1 => n3047, 
                           B2 => mult_143_n5626, C1 => mult_143_n5625, C2 => 
                           mult_143_n5626, ZN => mult_143_n5617);
   U1383 : INV_X1 port map( A => n4727, ZN => n4688);
   U1389 : AOI222_X1 port map( A1 => mult_143_n2759, A2 => mult_143_n6367, B1 
                           => mult_143_n2759, B2 => mult_143_n6368, C1 => 
                           mult_143_n6367, C2 => mult_143_n6368, ZN => n4689);
   U1392 : XNOR2_X1 port map( A => n3803, B => mult_143_n5953, ZN => n3116);
   U1393 : XOR2_X1 port map( A => mult_143_n4972, B => mult_143_n4973, Z => 
                           n4690);
   U1411 : OR2_X1 port map( A1 => mult_143_n5284, A2 => mult_143_n5285, ZN => 
                           n4772);
   U1439 : INV_X1 port map( A => n4693, ZN => n4694);
   U1442 : INV_X1 port map( A => n4748, ZN => n4695);
   U1444 : AOI222_X1 port map( A1 => n994, A2 => n970, B1 => n970, B2 => 
                           mult_143_n5662, C1 => mult_143_n5662, C2 => n994, ZN
                           => mult_143_n5650);
   U1448 : OAI21_X1 port map( B1 => mult_143_n6549, B2 => n3117, A => 
                           mult_143_n4767, ZN => mult_143_n4787);
   U1449 : XOR2_X1 port map( A => n419, B => mult_143_n5594, Z => 
                           mult_143_n5593);
   U1450 : XNOR2_X1 port map( A => mult_143_n5593, B => mult_143_n5631, ZN => 
                           mult_143_n5571);
   U1451 : XNOR2_X1 port map( A => n1749, B => mult_143_n5321, ZN => n4699);
   U1452 : XOR2_X1 port map( A => n4872, B => mult_143_n4852, Z => n4700);
   U1453 : XOR2_X1 port map( A => mult_143_n4948, B => mult_143_n4949, Z => 
                           n4701);
   U1475 : AOI222_X1 port map( A1 => n3108, A2 => n964, B1 => n3108, B2 => 
                           mult_143_n5670, C1 => n964, C2 => mult_143_n5670, ZN
                           => mult_143_n5656);
   U1476 : XNOR2_X1 port map( A => n4702, B => n4703, ZN => n1045);
   U1477 : XNOR2_X1 port map( A => n1677, B => n3698, ZN => n4703);
   U1478 : XNOR2_X1 port map( A => mult_143_n5345, B => n4704, ZN => 
                           mult_143_n5263);
   U1479 : XOR2_X1 port map( A => mult_143_n5346, B => mult_143_n5347, Z => 
                           n4704);
   U1485 : XNOR2_X1 port map( A => n3491, B => n3598, ZN => n4710);
   U1488 : AOI222_X1 port map( A1 => n1474, A2 => n1597, B1 => n4842, B2 => 
                           n3696, C1 => n1597, C2 => n3696, ZN => 
                           mult_143_n5446);
   U1489 : XNOR2_X1 port map( A => n4981, B => mult_143_n4989, ZN => n4713);
   U1490 : INV_X1 port map( A => n4743, ZN => n4714);
   U1491 : XNOR2_X1 port map( A => n1528, B => n4749, ZN => mult_143_n4984);
   U1492 : XNOR2_X1 port map( A => n4716, B => n4717, ZN => n1562);
   U1493 : XNOR2_X1 port map( A => n4718, B => n3830, ZN => mult_143_n5189);
   U1494 : XNOR2_X1 port map( A => n3706, B => n1562, ZN => n4718);
   U1495 : XNOR2_X1 port map( A => n3066, B => n4798, ZN => mult_143_n5743);
   U1496 : XNOR2_X1 port map( A => mult_143_n5669, B => n453, ZN => n4720);
   U1497 : OAI22_X1 port map( A1 => n3000, A2 => mult_143_n6421, B1 => n3093, 
                           B2 => n2711, ZN => mult_143_n5479);
   U1498 : XOR2_X1 port map( A => n4721, B => n3583, Z => n3091);
   U1499 : INV_X1 port map( A => n4722, ZN => n4723);
   U1506 : OR2_X1 port map( A1 => mult_143_n5578, A2 => n1478, ZN => n4724);
   U1508 : XNOR2_X1 port map( A => mult_143_n5739, B => n4725, ZN => n2770);
   U1510 : XNOR2_X1 port map( A => n3500, B => n3738, ZN => mult_143_n5414);
   U1511 : XOR2_X1 port map( A => n4699, B => n3726, Z => n4726);
   U1513 : INV_X1 port map( A => mult_143_n5352, ZN => n4781);
   U1514 : XNOR2_X1 port map( A => mult_143_n5254, B => mult_143_n5253, ZN => 
                           n387);
   U1515 : XNOR2_X1 port map( A => mult_143_n5351, B => n4781, ZN => 
                           mult_143_n5254);
   U1516 : CLKBUF_X1 port map( A => mult_143_n426, Z => n4728);
   U1518 : AOI222_X1 port map( A1 => n698, A2 => n4652, B1 => n698, B2 => n2664
                           , C1 => n4950, C2 => n2664, ZN => n4729);
   U1519 : XNOR2_X1 port map( A => n4730, B => n3584, ZN => n1651);
   U1520 : OAI22_X1 port map( A1 => n2847, A2 => n4792, B1 => mult_143_n6360, 
                           B2 => n2613, ZN => mult_143_n5730);
   U1521 : XNOR2_X1 port map( A => n4806, B => n1757, ZN => mult_143_n5276);
   U1524 : XNOR2_X1 port map( A => mult_143_n5341, B => mult_143_n5338, ZN => 
                           n4732);
   U1525 : INV_X1 port map( A => n4733, ZN => n4734);
   U1528 : OAI22_X1 port map( A1 => n4738, A2 => n4746, B1 => n4739, B2 => 
                           n4735, ZN => n4737);
   U1529 : XNOR2_X1 port map( A => mult_143_n5944, B => n3803, ZN => 
                           mult_143_n6401);
   U1532 : AOI21_X1 port map( B1 => mult_143_n4759, B2 => n2784, A => 
                           mult_143_n6560, ZN => n4742);
   U1533 : XNOR2_X1 port map( A => n2844, B => mult_143_n1690, ZN => 
                           mult_143_n5557);
   U1534 : AOI222_X1 port map( A1 => n740, A2 => n968, B1 => n968, B2 => 
                           mult_143_n5586, C1 => n740, C2 => mult_143_n5586, ZN
                           => n4744);
   U1535 : AOI222_X1 port map( A1 => n740, A2 => n968, B1 => n968, B2 => 
                           mult_143_n5586, C1 => n740, C2 => mult_143_n5586, ZN
                           => mult_143_n5612);
   U1536 : OAI22_X1 port map( A1 => n4782, A2 => mult_143_n5174, B1 => n991, B2
                           => n4949, ZN => mult_143_n5180);
   U1537 : NAND2_X1 port map( A1 => n4736, A2 => n3817, ZN => n4778);
   U1538 : AND2_X1 port map( A1 => n4949, A2 => n991, ZN => n4782);
   U1541 : XOR2_X1 port map( A => n4749, B => n4751, Z => n1621);
   U1542 : OAI22_X1 port map( A1 => mult_143_n5163, A2 => n4794, B1 => 
                           mult_143_n5164, B2 => n3105, ZN => n2909);
   U1543 : XNOR2_X1 port map( A => n1045, B => n1050, ZN => mult_143_n5568);
   U1545 : XNOR2_X1 port map( A => mult_143_n5016, B => n4752, ZN => n1629);
   U1548 : OAI21_X1 port map( B1 => mult_143_n4340, B2 => mult_143_n4784, A => 
                           mult_143_n4475, ZN => n4756);
   U1549 : OAI222_X1 port map( A1 => n4627, A2 => n4614, B1 => n4627, B2 => 
                           n4655, C1 => n4614, C2 => n4655, ZN => n2938);
   U1551 : XNOR2_X1 port map( A => mult_143_n5568, B => n1066, ZN => n4758);
   U1552 : OAI22_X1 port map( A1 => n4799, A2 => n4754, B1 => n3066, B2 => 
                           n4638, ZN => mult_143_n5765);
   U1553 : INV_X1 port map( A => n3797, ZN => n1839);
   U1557 : XNOR2_X1 port map( A => n4784, B => n3768, ZN => n1042);
   U1558 : AOI222_X1 port map( A1 => n3671, A2 => n3732, B1 => n3671, B2 => 
                           n3492, C1 => n3495, C2 => n3732, ZN => n4762);
   U1559 : XNOR2_X1 port map( A => mult_143_n5682, B => n3734, ZN => n4763);
   U1561 : AOI222_X1 port map( A1 => n3671, A2 => n3732, B1 => n3671, B2 => 
                           n3492, C1 => n3495, C2 => n4853, ZN => n1471);
   U1562 : NOR2_X1 port map( A1 => n4817, A2 => n4816, ZN => n4815);
   U1563 : AOI222_X1 port map( A1 => n4874, A2 => mult_143_n5616, B1 => n4874, 
                           B2 => n4875, C1 => n4875, C2 => mult_143_n5616, ZN 
                           => n4764);
   U1565 : XNOR2_X1 port map( A => n2938, B => n3636, ZN => n4806);
   U1567 : XNOR2_X1 port map( A => n4776, B => n4760, ZN => n3066);
   U1568 : BUF_X2 port map( A => n3790, Z => n4765);
   U1569 : AOI222_X1 port map( A1 => n2739, A2 => mult_143_n6367, B1 => n2739, 
                           B2 => n4602, C1 => n4670, C2 => n4602, ZN => 
                           mult_143_n5422);
   U1572 : XNOR2_X1 port map( A => n4807, B => n2840, ZN => n3051);
   U1573 : NAND2_X1 port map( A1 => n3775, A2 => n4747, ZN => mult_143_n1898);
   U1574 : NAND2_X1 port map( A1 => n3775, A2 => n4845, ZN => mult_143_n1902);
   U1575 : NAND2_X1 port map( A1 => n3775, A2 => n4736, ZN => mult_143_n1900);
   U1576 : XOR2_X1 port map( A => n4770, B => n4771, Z => n4769);
   U1578 : NAND4_X1 port map( A1 => n4773, A2 => n1008, A3 => n4772, A4 => 
                           n4600, ZN => n584);
   U1579 : INV_X1 port map( A => n2875, ZN => n4773);
   U1580 : NOR2_X1 port map( A1 => n2850, A2 => n961, ZN => n4774);
   U1581 : AOI21_X1 port map( B1 => n2850, B2 => n961, A => mult_143_n5422, ZN 
                           => n4775);
   U1582 : NAND2_X1 port map( A1 => n3020, A2 => n3071, ZN => n4776);
   U1583 : NOR2_X1 port map( A1 => n4779, A2 => n4777, ZN => n1536);
   U1584 : OAI21_X1 port map( B1 => n3675, B2 => n3673, A => n4778, ZN => n4777
                           );
   U1585 : INV_X1 port map( A => mult_143_n5943, ZN => n4779);
   U1586 : XNOR2_X1 port map( A => n4886, B => mult_143_n5556, ZN => n3118);
   U1588 : XNOR2_X1 port map( A => n3729, B => n1669, ZN => n4780);
   U1589 : OAI22_X1 port map( A1 => n1691, A2 => n4820, B1 => n3682, B2 => 
                           n3723, ZN => mult_143_n1005);
   U1590 : XNOR2_X1 port map( A => mult_143_n4919, B => n4754, ZN => 
                           mult_143_n4915);
   U1591 : XNOR2_X1 port map( A => n2739, B => n4730, ZN => mult_143_n5610);
   U1593 : NAND2_X1 port map( A1 => n4787, A2 => n4786, ZN => mult_143_n5080);
   U1594 : AOI22_X1 port map( A1 => n4631, A2 => n4626, B1 => n3784, B2 => 
                           n3531, ZN => n4786);
   U1595 : NAND2_X1 port map( A1 => n4695, A2 => n3820, ZN => n4787);
   U1596 : INV_X1 port map( A => mult_143_n6346, ZN => n4789);
   U1597 : AOI21_X1 port map( B1 => n4688, B2 => n3820, A => n4813, ZN => n4812
                           );
   U1598 : AND2_X1 port map( A1 => n3106, A2 => mult_143_n5164, ZN => n4790);
   U1599 : OAI22_X1 port map( A1 => n4791, A2 => mult_143_n5378, B1 => 
                           mult_143_n5377, B2 => n4686, ZN => n1484);
   U1600 : AND2_X1 port map( A1 => mult_143_n5376, A2 => mult_143_n5377, ZN => 
                           n4791);
   U1601 : AOI21_X1 port map( B1 => n4769, B2 => n4589, A => n2765, ZN => n2953
                           );
   U1602 : AND2_X1 port map( A1 => n2613, A2 => mult_143_n6360, ZN => n4792);
   U1603 : XNOR2_X1 port map( A => n2621, B => n4793, ZN => mult_143_n5273);
   U1604 : XNOR2_X1 port map( A => n2728, B => mult_143_n5363, ZN => n4793);
   U1605 : XNOR2_X1 port map( A => n1627, B => n4624, ZN => mult_143_n4928);
   U1607 : AND2_X1 port map( A1 => n3105, A2 => mult_143_n5164, ZN => n4794);
   U1608 : XNOR2_X1 port map( A => n3054, B => mult_143_n1896, ZN => n4795);
   U1609 : OAI21_X1 port map( B1 => n4797, B2 => n4796, A => n4574, ZN => n1490
                           );
   U1610 : AND2_X1 port map( A1 => mult_143_n5505, A2 => mult_143_n5508, ZN => 
                           n4796);
   U1611 : INV_X1 port map( A => mult_143_n5507, ZN => n4797);
   U1612 : AND2_X1 port map( A1 => n3066, A2 => n4638, ZN => n4799);
   U1613 : XNOR2_X1 port map( A => n4673, B => n4800, ZN => mult_143_n5769);
   U1614 : INV_X1 port map( A => mult_143_n5760, ZN => n4800);
   U1615 : NAND2_X1 port map( A1 => n4805, A2 => n4802, ZN => mult_143_n4920);
   U1616 : INV_X1 port map( A => n4803, ZN => n4802);
   U1617 : OAI21_X1 port map( B1 => n3644, B2 => n3613, A => n4804, ZN => n4803
                           );
   U1618 : NAND2_X1 port map( A1 => n4695, A2 => n3538, ZN => n4804);
   U1619 : NAND2_X1 port map( A1 => n4688, A2 => n3807, ZN => n4805);
   U1620 : OAI21_X1 port map( B1 => n3050, B2 => n4810, A => n4635, ZN => n4809
                           );
   U1621 : AND2_X1 port map( A1 => n2726, A2 => n3795, ZN => n4810);
   U1622 : INV_X1 port map( A => mult_143_n652, ZN => mult_143_n4510);
   U1623 : AND2_X1 port map( A1 => mult_143_n652, A2 => n4811, ZN => 
                           mult_143_n5528);
   U1624 : NAND2_X1 port map( A1 => mult_143_n6581, A2 => mult_143_n6582, ZN =>
                           n4811);
   U1625 : NAND2_X1 port map( A1 => n4814, A2 => n4812, ZN => mult_143_n5090);
   U1626 : NOR2_X1 port map( A1 => n3643, A2 => n3613, ZN => n4813);
   U1627 : NAND2_X1 port map( A1 => n4695, A2 => n3531, ZN => n4814);
   U1628 : XNOR2_X1 port map( A => n4815, B => mult_143_n5166, ZN => 
                           mult_143_n5417);
   U1629 : NOR2_X1 port map( A1 => mult_143_n5419, A2 => mult_143_n6381, ZN => 
                           n4816);
   U1630 : AOI21_X1 port map( B1 => mult_143_n5419, B2 => mult_143_n6381, A => 
                           mult_143_n5420, ZN => n4817);
   U1631 : OAI22_X1 port map( A1 => n4819, A2 => n4818, B1 => mult_143_n5481, 
                           B2 => n4674, ZN => n1489);
   U1632 : INV_X1 port map( A => mult_143_n5483, ZN => n4818);
   U1633 : AND2_X1 port map( A1 => n3682, A2 => n3723, ZN => n4820);
   U1634 : XNOR2_X1 port map( A => mult_143_n6365, B => n4753, ZN => n4821);
   U1635 : NAND2_X1 port map( A1 => n3531, A2 => n4766, ZN => mult_143_n1942);
   U1636 : NAND2_X1 port map( A1 => n2840, A2 => n4688, ZN => mult_143_n1895);
   MY_CLK_r_REG1379_S1 : DFF_X1 port map( D => n1610, CK => clk, Q => n_1390, 
                           QN => n4621);
   MY_CLK_r_REG1177_S2 : DFF_X1 port map( D => n606, CK => clk, Q => n_1391, QN
                           => n4717);
   MY_CLK_r_REG1182_S2 : DFF_X1 port map( D => mult_143_n5702, CK => clk, Q => 
                           n4926, QN => n4568);
   U1185 : XNOR2_X2 port map( A => mult_143_n6270, B => B_SIG(7), ZN => 
                           mult_143_n2798);
   MY_CLK_r_REG1159_S2 : DFF_X1 port map( D => n1693, CK => clk, Q => n3738, QN
                           => n_1392);
   MY_CLK_r_REG1373_S1 : DFF_X1 port map( D => mult_143_n6621, CK => clk, Q => 
                           n3539, QN => n4719);
   MY_CLK_r_REG1500_S1 : DFF_X1 port map( D => B_SIG(12), CK => clk, Q => n3779
                           , QN => n4667);
   MY_CLK_r_REG1148_S2 : DFF_X1 port map( D => n1477, CK => clk, Q => n3500, QN
                           => n_1393);
   MY_CLK_r_REG1466_S1 : DFF_X2 port map( D => n1030, CK => clk, Q => n3771, QN
                           => n4693);
   MY_CLK_r_REG1189_S2 : DFF_X1 port map( D => n2945, CK => clk, Q => n3491, QN
                           => n4861);
   MY_CLK_r_REG1199_S2 : DFF_X1 port map( D => n1482, CK => clk, Q => n3506, QN
                           => n4868);
   U1554 : NAND2_X1 port map( A1 => n3782, A2 => n3809, ZN => n4785);
   U170 : XNOR2_X1 port map( A => B_SIG(3), B => mult_143_n6230, ZN => 
                           mult_143_n6630);
   U1484 : INV_X1 port map( A => mult_143_n3083, ZN => n4709);
   MY_CLK_r_REG1211_S2 : DFF_X1 port map( D => n1469, CK => clk, Q => n3493, QN
                           => n_1394);
   MY_CLK_r_REG1487_S1 : DFF_X1 port map( D => B_SIG(17), CK => clk, Q => n3784
                           , QN => n4889);
   MY_CLK_r_REG1443_S1 : DFF_X1 port map( D => n1026, CK => clk, Q => n3808, QN
                           => n_1395);
   U6 : OR2_X1 port map( A1 => n2688, A2 => n3099, ZN => n2666);
   U78 : AOI22_X1 port map( A1 => n734, A2 => mult_143_n6551, B1 => n972, B2 =>
                           mult_143_n5677, ZN => n4833);
   U126 : XNOR2_X1 port map( A => n3139, B => n3099, ZN => n3047);
   U176 : AOI222_X1 port map( A1 => mult_143_n6479, A2 => mult_143_n6478, B1 =>
                           mult_143_n6478, B2 => n4583, C1 => mult_143_n6479, 
                           C2 => n4583, ZN => mult_143_n5350);
   U210 : OR2_X1 port map( A1 => mult_143_n5143, A2 => mult_143_n5144, ZN => 
                           n4901);
   U220 : XNOR2_X1 port map( A => mult_143_n5844, B => mult_143_n6367, ZN => 
                           n3090);
   U234 : INV_X1 port map( A => mult_143_n3154, ZN => n4860);
   U247 : AND2_X1 port map( A1 => n3506, A2 => n3728, ZN => n4831);
   U280 : AND2_X1 port map( A1 => n3801, A2 => n3827, ZN => n4835);
   U296 : NOR2_X1 port map( A1 => mult_143_n5815, A2 => n4835, ZN => 
                           mult_143_n5814);
   U310 : AND2_X1 port map( A1 => n3800, A2 => n3820, ZN => n4834);
   U331 : XNOR2_X1 port map( A => n4880, B => n4830, ZN => n1633);
   U371 : OAI21_X1 port map( B1 => B_SIG(3), B2 => B_SIG(1), A => B_SIG(2), ZN 
                           => mult_143_n6308);
   U386 : INV_X1 port map( A => n4889, ZN => n4890);
   U391 : OR2_X1 port map( A1 => mult_143_n5169, A2 => mult_143_n5168, ZN => 
                           n2936);
   U425 : INV_X1 port map( A => B_SIG(3), ZN => n909);
   U516 : INV_X1 port map( A => n4750, ZN => n2751);
   U575 : INV_X1 port map( A => mult_143_n5676, ZN => n4832);
   U707 : INV_X1 port map( A => B_SIG(0), ZN => n629);
   U725 : NAND2_X1 port map( A1 => n2881, A2 => mult_143_n5261, ZN => 
                           mult_143_n5260);
   U843 : AOI222_X1 port map( A1 => mult_143_n6361, A2 => mult_143_n6362, B1 =>
                           mult_143_n6361, B2 => n2704, C1 => mult_143_n6362, 
                           C2 => n2704, ZN => mult_143_n5718);
   U852 : CLKBUF_X1 port map( A => mult_143_n3239, Z => n1030);
   U853 : OR2_X1 port map( A1 => n3506, A2 => n3728, ZN => n4827);
   U873 : AND2_X1 port map( A1 => mult_143_n5242, A2 => n1037, ZN => n4828);
   U945 : INV_X1 port map( A => n4879, ZN => n4830);
   U951 : OAI21_X1 port map( B1 => n4831, B2 => n1675, A => n4827, ZN => n2911)
                           ;
   U999 : XNOR2_X1 port map( A => n4833, B => n4832, ZN => n1644);
   U1001 : NOR2_X1 port map( A1 => mult_143_n5017, A2 => n4834, ZN => 
                           mult_143_n5016);
   U1002 : OAI211_X1 port map( C1 => n3655, C2 => n3597, A => n4785, B => 
                           mult_143_n5892, ZN => n4784);
   U1006 : OAI22_X1 port map( A1 => n4836, A2 => mult_143_n5477, B1 => 
                           mult_143_n5478, B2 => mult_143_n5479, ZN => 
                           mult_143_n5483);
   U1030 : AND2_X1 port map( A1 => mult_143_n5479, A2 => mult_143_n5478, ZN => 
                           n4836);
   U1043 : XNOR2_X1 port map( A => n1749, B => n4837, ZN => n2885);
   U1057 : XNOR2_X1 port map( A => mult_143_n5321, B => n3726, ZN => n4837);
   U1062 : XNOR2_X1 port map( A => mult_143_n5664, B => mult_143_n6513, ZN => 
                           mult_143_n5182);
   U1067 : OAI22_X1 port map( A1 => n1574, A2 => n4657, B1 => n2685, B2 => 
                           n4625, ZN => n4838);
   U1073 : XNOR2_X1 port map( A => mult_143_n5772, B => mult_143_n4490, ZN => 
                           n4839);
   U1096 : XNOR2_X1 port map( A => n4759, B => n1542, ZN => n2750);
   U1104 : XOR2_X1 port map( A => mult_143_n5667, B => mult_143_n5668, Z => 
                           n4841);
   U1135 : AOI222_X1 port map( A1 => n3610, A2 => n3829, B1 => n3610, B2 => 
                           n3499, C1 => n3829, C2 => n3499, ZN => n4842);
   U1155 : OAI222_X1 port map( A1 => n4933, A2 => n4581, B1 => n4933, B2 => 
                           n4582, C1 => n4581, C2 => n4582, ZN => n4843);
   U1160 : XNOR2_X1 port map( A => n4754, B => mult_143_n1610, ZN => 
                           mult_143_n5751);
   U1161 : XNOR2_X1 port map( A => n1563, B => n3793, ZN => mult_143_n4973);
   U1173 : XNOR2_X1 port map( A => mult_143_n5354, B => n4844, ZN => 
                           mult_143_n5266);
   U1179 : XNOR2_X1 port map( A => mult_143_n5355, B => mult_143_n5356, ZN => 
                           n4844);
   U1194 : INV_X1 port map( A => n4667, ZN => n4845);
   U1219 : XNOR2_X1 port map( A => mult_143_n5728, B => n4847, ZN => n4859);
   U1221 : XOR2_X1 port map( A => mult_143_n4504, B => mult_143_n5751, Z => 
                           n4847);
   U1222 : INV_X1 port map( A => n4680, ZN => n4848);
   U1227 : XNOR2_X1 port map( A => n4849, B => n4850, ZN => n1561);
   U1249 : NOR2_X1 port map( A1 => n3488, A2 => n3608, ZN => n4928);
   U1257 : OR2_X1 port map( A1 => n3594, A2 => n3613, ZN => n4921);
   U1270 : OAI211_X1 port map( C1 => n3527, C2 => n3554, A => n3668, B => n3601
                           , ZN => n4851);
   U1290 : AND2_X1 port map( A1 => n3539, A2 => n3778, ZN => n4912);
   U1301 : AND2_X1 port map( A1 => n4932, A2 => n4930, ZN => n4755);
   U1306 : INV_X1 port map( A => n4852, ZN => n4853);
   U1326 : XNOR2_X1 port map( A => n4854, B => n4855, ZN => n3027);
   U1371 : CLKBUF_X1 port map( A => mult_143_n2702, Z => n4856);
   U1480 : AOI222_X1 port map( A1 => n972, A2 => mult_143_n5676, B1 => 
                           mult_143_n5677, B2 => n972, C1 => mult_143_n5677, C2
                           => mult_143_n5676, ZN => n4857);
   U1481 : AOI222_X1 port map( A1 => n972, A2 => mult_143_n5676, B1 => 
                           mult_143_n5677, B2 => n972, C1 => mult_143_n5677, C2
                           => mult_143_n5676, ZN => mult_143_n5688);
   U1483 : XNOR2_X1 port map( A => mult_143_n4504, B => mult_143_n5751, ZN => 
                           n4858);
   U1486 : XNOR2_X1 port map( A => n4859, B => mult_143_n5725, ZN => n1646);
   U1522 : XNOR2_X1 port map( A => n4861, B => n4862, ZN => n1683);
   U1531 : XNOR2_X1 port map( A => mult_143_n5854, B => n3791, ZN => n4863);
   U1544 : XNOR2_X1 port map( A => mult_143_n5570, B => mult_143_n5569, ZN => 
                           n4864);
   U1547 : XNOR2_X1 port map( A => n4826, B => n3731, ZN => n1631);
   U1570 : NOR2_X1 port map( A1 => n4866, A2 => n4867, ZN => n1008);
   U1637 : AND2_X1 port map( A1 => n2934, A2 => n542, ZN => n4866);
   U1638 : NOR2_X1 port map( A1 => n4726, A2 => mult_143_n5285, ZN => n4867);
   U1639 : XOR2_X1 port map( A => n4868, B => n4869, Z => n4883);
   U1640 : XNOR2_X1 port map( A => n3703, B => n3505, ZN => n1675);
   U1641 : OAI21_X1 port map( B1 => n605, B2 => mult_143_n4502, A => n604, ZN 
                           => n4870);
   U1642 : INV_X1 port map( A => n4743, ZN => n4871);
   U1643 : OR2_X1 port map( A1 => n4929, A2 => n4928, ZN => n4927);
   U1644 : NAND2_X1 port map( A1 => n1678, A2 => n4927, ZN => mult_143_n427);
   U1645 : XOR2_X1 port map( A => n1590, B => n1614, Z => n4872);
   U1646 : XNOR2_X1 port map( A => n4873, B => n2847, ZN => mult_143_n5722);
   U1647 : XNOR2_X1 port map( A => n2613, B => mult_143_n6360, ZN => n4873);
   U1648 : XOR2_X1 port map( A => mult_143_n5628, B => mult_143_n5619, Z => 
                           n4874);
   U1649 : AOI222_X1 port map( A1 => n3047, A2 => mult_143_n5625, B1 => n3047, 
                           B2 => mult_143_n5626, C1 => mult_143_n5625, C2 => 
                           mult_143_n5626, ZN => n4875);
   U1650 : NOR2_X2 port map( A1 => mult_143_n5637, A2 => n2768, ZN => 
                           mult_143_n5626);
   U1651 : AOI222_X4 port map( A1 => mult_143_n5345, A2 => mult_143_n5346, B1 
                           => mult_143_n5345, B2 => mult_143_n5347, C1 => 
                           mult_143_n5346, C2 => mult_143_n5347, ZN => 
                           mult_143_n5261);
   U1653 : XNOR2_X1 port map( A => n3660, B => n3745, ZN => n4877);
   U1654 : XOR2_X1 port map( A => n1629, B => mult_143_n5015, Z => n4878);
   U1656 : BUF_X1 port map( A => mult_143_n5204, Z => n4882);
   U1657 : INV_X2 port map( A => n4730, ZN => mult_143_n6367);
   U1658 : XNOR2_X1 port map( A => n1675, B => n4883, ZN => mult_143_n5607);
   U1660 : AOI222_X1 port map( A1 => n1648, A2 => n3555, B1 => n3555, B2 => 
                           n3737, C1 => n1648, C2 => n3737, ZN => n4885);
   U1661 : XNOR2_X1 port map( A => n2844, B => mult_143_n1690, ZN => n4886);
   U1662 : NAND2_X1 port map( A1 => mult_143_n5607, A2 => mult_143_n5606, ZN =>
                           n4887);
   U1663 : XNOR2_X1 port map( A => n2852, B => mult_143_n5422, ZN => n4888);
   U1665 : AOI21_X1 port map( B1 => n4870, B2 => n1056, A => mult_143_n335, ZN 
                           => n4892);
   U1667 : XNOR2_X1 port map( A => n4894, B => n4768, ZN => n1669);
   U1668 : XNOR2_X1 port map( A => n4895, B => n4896, ZN => n1559);
   U1670 : INV_X2 port map( A => n4759, ZN => n4760);
   U1674 : AND2_X1 port map( A1 => n3548, A2 => n3756, ZN => n4907);
   U1675 : OAI22_X1 port map( A1 => n1561, A2 => n4907, B1 => n3756, B2 => 
                           n3548, ZN => mult_143_n5606);
   U1676 : INV_X1 port map( A => n4901, ZN => mult_143_n6577);
   U1677 : OAI21_X1 port map( B1 => n4723, B2 => n3701, A => n3488, ZN => n4932
                           );
   U1678 : AOI21_X1 port map( B1 => n3488, B2 => n4723, A => n3701, ZN => n4929
                           );
   U1679 : AND2_X1 port map( A1 => n3728, A2 => n3506, ZN => n4909);
   U1680 : OAI22_X1 port map( A1 => n1675, A2 => n4909, B1 => n3728, B2 => 
                           n3506, ZN => mult_143_n5208);
   U1683 : XNOR2_X1 port map( A => n4903, B => n4904, ZN => n1578);
   U1685 : OAI22_X1 port map( A1 => n1631, A2 => n4908, B1 => n3752, B2 => 
                           n3513, ZN => mult_143_n5152);
   U1686 : AND2_X1 port map( A1 => n3752, A2 => n3513, ZN => n4908);
   U1687 : NAND2_X1 port map( A1 => mult_143_n5621, A2 => mult_143_n5601, ZN =>
                           n4910);
   U1689 : NOR2_X1 port map( A1 => mult_143_n5493, A2 => n4912, ZN => 
                           mult_143_n5492);
   U1697 : XNOR2_X1 port map( A => n3027, B => n4920, ZN => mult_143_n5739);
   U1698 : XNOR2_X1 port map( A => n3499, B => n4609, ZN => n4920);
   U1699 : NAND2_X1 port map( A1 => mult_143_n4981, A2 => n4921, ZN => 
                           mult_143_n4980);
   U1700 : NAND2_X1 port map( A1 => mult_143_n5374, A2 => mult_143_n5375, ZN =>
                           n3084);
   U1701 : XNOR2_X1 port map( A => n2905, B => mult_143_n5477, ZN => 
                           mult_143_n5374);
   U1702 : AOI21_X1 port map( B1 => n1042, B2 => n496, A => n4922, ZN => n3000)
                           ;
   U1703 : NAND2_X1 port map( A1 => n4923, A2 => n2711, ZN => n4922);
   U1704 : NAND2_X1 port map( A1 => n1657, A2 => n986, ZN => n4923);
   U1705 : NAND2_X1 port map( A1 => n4924, A2 => n4828, ZN => mult_143_n6619);
   U1706 : NAND3_X1 port map( A1 => n505, A2 => n516, A3 => n519, ZN => n4924);
   U1707 : NOR2_X2 port map( A1 => mult_143_n4809, A2 => mult_143_n5204, ZN => 
                           n1056);
   U1708 : XNOR2_X1 port map( A => n1687, B => n4925, ZN => mult_143_n5206);
   U1709 : XNOR2_X1 port map( A => n3735, B => n4926, ZN => n4925);
   U1710 : NAND2_X1 port map( A1 => n3608, A2 => n3701, ZN => n4930);
   MY_CLK_r_REG1238_S2 : DFF_X1 port map( D => n1702, CK => clk, Q => n3747, QN
                           => n_1396);
   MY_CLK_r_REG1146_S2 : DFF_X1 port map( D => n1710, CK => clk, Q => n3756, QN
                           => n4880);
   MY_CLK_r_REG1357_S2 : DFF_X1 port map( D => mult_143_n5256, CK => clk, Q => 
                           n3527, QN => n_1397);
   MY_CLK_r_REG1375_S1 : DFF_X1 port map( D => mult_143_n4820, CK => clk, Q => 
                           n3594, QN => n4589);
   MY_CLK_r_REG1378_S1 : DFF_X1 port map( D => n804, CK => clk, Q => n3767, QN 
                           => n_1398);
   MY_CLK_r_REG1376_S1 : DFF_X1 port map( D => n649, CK => clk, Q => n3773, QN 
                           => n4632);
   MY_CLK_r_REG1429_S1 : DFF_X1 port map( D => A_SIG(5), CK => clk, Q => n3792,
                           QN => n4590);
   MY_CLK_r_REG1401_S1 : DFF_X1 port map( D => mult_143_n4828, CK => clk, Q => 
                           n3644, QN => n4733);
   MY_CLK_r_REG1454_S1 : DFF_X1 port map( D => mult_143_n5124, CK => clk, Q => 
                           n3659, QN => n_1399);
   U437 : INV_X1 port map( A => n4749, ZN => n4750);
   U1555 : INV_X1 port map( A => n3768, ZN => n2864);
   U414 : INV_X1 port map( A => n4721, ZN => n3099);
   U225 : INV_X1 port map( A => n3796, ZN => n2780);
   U1682 : OAI22_X1 port map( A1 => n2794, A2 => n3120, B1 => n3510, B2 => 
                           n3742, ZN => n2890);
   U510 : AOI222_X1 port map( A1 => n2874, A2 => n2829, B1 => n2874, B2 => 
                           n3057, C1 => n2829, C2 => n3057, ZN => 
                           mult_143_n5586);
   U466 : OAI21_X1 port map( B1 => mult_143_n4788, B2 => mult_143_n4789, A => 
                           mult_143_n6550, ZN => mult_143_n4766);
   U16 : INV_X1 port map( A => B_SIG(1), ZN => n630);
   U416 : NAND2_X1 port map( A1 => B_SIG(1), A2 => B_SIG(0), ZN => 
                           mult_143_n6296);
   MY_CLK_r_REG1364_S1 : DFF_X1 port map( D => n2599, CK => clk, Q => n3805, QN
                           => n4692);
   MY_CLK_r_REG1140_S2 : DFF_X1 port map( D => n1480, CK => clk, Q => n3503, QN
                           => n4571);
   MY_CLK_r_REG1193_S2 : DFF_X1 port map( D => n1644, CK => clk, Q => n3706, QN
                           => n_1400);
   MY_CLK_r_REG1170_S2 : DFF_X1 port map( D => n1472, CK => clk, Q => n3497, QN
                           => n4876);
   MY_CLK_r_REG1393_S1 : DFF_X1 port map( D => n765, CK => clk, Q => n3802, QN 
                           => n4680);
   MY_CLK_r_REG1214_S2 : DFF_X1 port map( D => n1475, CK => clk, Q => n3498, QN
                           => n_1401);
   U8 : CLKBUF_X1 port map( A => mult_143_n427, Z => n4731);
   U25 : AOI222_X1 port map( A1 => mult_143_n6417, A2 => n4575, B1 => 
                           mult_143_n6417, B2 => n2622, C1 => n4575, C2 => 
                           n2622, ZN => mult_143_n5556);
   U29 : AOI222_X1 port map( A1 => mult_143_n6590, A2 => n1628, B1 => 
                           mult_143_n6590, B2 => mult_143_n6592, C1 => n1628, 
                           C2 => mult_143_n6592, ZN => mult_143_n5676);
   U30 : AOI222_X1 port map( A1 => mult_143_n5333, A2 => n2725, B1 => 
                           mult_143_n5334, B2 => mult_143_n5333, C1 => 
                           mult_143_n5334, C2 => n2725, ZN => mult_143_n5322);
   U31 : OAI22_X1 port map( A1 => n4937, A2 => mult_143_n6589, B1 => 
                           mult_143_n4989, B2 => n4981, ZN => mult_143_n5677);
   U41 : OR2_X1 port map( A1 => n2994, A2 => n2993, ZN => mult_143_n5381);
   U61 : NAND2_X1 port map( A1 => mult_143_n5578, A2 => n1478, ZN => 
                           mult_143_n412);
   U73 : NAND2_X1 port map( A1 => n4968, A2 => n4967, ZN => n1478);
   U74 : NAND2_X1 port map( A1 => n4970, A2 => n4969, ZN => n4968);
   U96 : AND2_X1 port map( A1 => n3802, A2 => n4675, ZN => n4979);
   U221 : INV_X1 port map( A => n1664, ZN => n4933);
   U338 : INV_X1 port map( A => mult_143_n5640, ZN => n4945);
   U375 : NAND2_X1 port map( A1 => n4945, A2 => n4944, ZN => n4943);
   U380 : AND2_X1 port map( A1 => n4766, A2 => n3801, ZN => n4966);
   U392 : NAND2_X1 port map( A1 => n3749, A2 => n3592, ZN => n4970);
   U401 : AND2_X1 port map( A1 => n3802, A2 => n3780, ZN => n4965);
   U445 : AND2_X1 port map( A1 => n3789, A2 => n3802, ZN => n4971);
   U479 : OR2_X1 port map( A1 => n3749, A2 => n3669, ZN => n4967);
   U513 : NOR2_X1 port map( A1 => mult_143_n5972, A2 => n4965, ZN => n3097);
   U520 : NOR2_X1 port map( A1 => mult_143_n5975, A2 => n4979, ZN => 
                           mult_143_n5974);
   U553 : INV_X1 port map( A => n4746, ZN => n4747);
   U556 : NOR2_X1 port map( A1 => mult_143_n5984, A2 => n4971, ZN => n1502);
   U637 : XNOR2_X1 port map( A => n4877, B => n4876, ZN => mult_143_n5639);
   U650 : AOI222_X1 port map( A1 => n3091, A2 => n4587, B1 => n3091, B2 => 
                           n2865, C1 => n4587, C2 => n2865, ZN => 
                           mult_143_n5341);
   U755 : AND2_X1 port map( A1 => n4981, A2 => mult_143_n4989, ZN => n4937);
   U822 : AND2_X1 port map( A1 => mult_143_n6555, A2 => n2717, ZN => n3030);
   U840 : AOI222_X1 port map( A1 => mult_143_n6382, A2 => n3116, B1 => 
                           mult_143_n6382, B2 => n4607, C1 => n3116, C2 => 
                           n4607, ZN => n2850);
   U1016 : INV_X1 port map( A => B_SIG(2), ZN => n910);
   U1094 : INV_X1 port map( A => n3774, ZN => n2895);
   U1146 : INV_X1 port map( A => n4753, ZN => n4754);
   U1152 : NAND2_X1 port map( A1 => n4939, A2 => n4938, ZN => mult_143_n6555);
   U1156 : OAI22_X1 port map( A1 => n3030, A2 => mult_143_n6554, B1 => 
                           mult_143_n6555, B2 => n2717, ZN => mult_143_n5719);
   U1243 : OAI21_X1 port map( B1 => B_SIG(1), B2 => B_SIG(0), A => 
                           mult_143_n6296, ZN => mult_143_n2458);
   U1327 : CLKBUF_X1 port map( A => mult_143_n4787, Z => n4697);
   U1482 : XOR2_X1 port map( A => n1617, B => mult_143_n4815, Z => n4935);
   U1539 : OR3_X1 port map( A1 => mult_143_n5639, A2 => mult_143_n5640, A3 => 
                           n4940, ZN => n4936);
   U1550 : NAND2_X1 port map( A1 => n2688, A2 => n3099, ZN => n4938);
   U1560 : NAND2_X1 port map( A1 => n1568, A2 => n3792, ZN => n4939);
   U1566 : AND2_X1 port map( A1 => n4636, A2 => n4829, ZN => n4940);
   U1571 : OAI211_X1 port map( C1 => n3643, C2 => n3675, A => n4942, B => n4941
                           , ZN => mult_143_n5033);
   U1606 : NAND2_X1 port map( A1 => n3772, A2 => n3782, ZN => n4941);
   U1652 : NAND2_X1 port map( A1 => n4736, A2 => n3820, ZN => n4942);
   U1671 : NOR2_X1 port map( A1 => n4943, A2 => mult_143_n5639, ZN => n4663);
   U1672 : NAND2_X1 port map( A1 => n4636, A2 => n4829, ZN => n4944);
   U1681 : XNOR2_X1 port map( A => n3572, B => n4590, ZN => n1664);
   U1684 : OAI22_X1 port map( A1 => mult_143_n5667, A2 => n546, B1 => n3678, B2
                           => n971, ZN => n4946);
   U1692 : OAI21_X1 port map( B1 => mult_143_n5656, B2 => n3038, A => n3036, ZN
                           => n4947);
   U1693 : NAND2_X1 port map( A1 => n4980, A2 => n4910, ZN => n740);
   U1695 : OAI21_X1 port map( B1 => n3130, B2 => mult_143_n4915, A => n4569, ZN
                           => n4949);
   U1711 : XOR2_X1 port map( A => mult_143_n5087, B => mult_143_n5086, Z => 
                           n4950);
   U1712 : XNOR2_X1 port map( A => mult_143_n5254, B => mult_143_n5253, ZN => 
                           n4951);
   U1713 : XNOR2_X1 port map( A => mult_143_n4510, B => n4952, ZN => 
                           mult_143_n5515);
   U1714 : XOR2_X1 port map( A => mult_143_n6581, B => mult_143_n6582, Z => 
                           n4952);
   U1716 : OAI22_X1 port map( A1 => mult_143_n5324, A2 => mult_143_n5325, B1 =>
                           mult_143_n5322, B2 => mult_143_n5323, ZN => n4955);
   U1717 : XNOR2_X1 port map( A => n4632, B => n4956, ZN => n1691);
   U1722 : XNOR2_X1 port map( A => n1507, B => n4721, ZN => mult_143_n1753);
   U1723 : XNOR2_X1 port map( A => n4963, B => n4964, ZN => n1597);
   U1724 : NOR2_X1 port map( A1 => n1525, A2 => n4966, ZN => mult_143_n5850);
   U1725 : INV_X1 port map( A => n3489, ZN => n4969);
   U1726 : OAI22_X1 port map( A1 => n4973, A2 => n4972, B1 => mult_143_n5654, 
                           B2 => mult_143_n5653, ZN => n1472);
   U1727 : OAI22_X1 port map( A1 => n4801, A2 => mult_143_n5180, B1 => 
                           mult_143_n5182, B2 => mult_143_n5181, ZN => n4972);
   U1728 : AND2_X1 port map( A1 => mult_143_n5653, A2 => mult_143_n5654, ZN => 
                           n4973);
   U1729 : OAI22_X1 port map( A1 => n1615, A2 => n3508, B1 => n3609, B2 => 
                           n3507, ZN => mult_143_n5240);
   U1730 : XNOR2_X1 port map( A => n4905, B => n4906, ZN => n1615);
   add_1_root_add_135_2 : FPmul_stage2_DW01_add_0 port map( A(7) => A_EXP(7), 
                           A(6) => A_EXP(6), A(5) => A_EXP(5), A(4) => A_EXP(4)
                           , A(3) => A_EXP(3), A(2) => A_EXP(2), A(1) => 
                           A_EXP(1), A(0) => A_EXP(0), B(7) => B_EXP(7), B(6) 
                           => B_EXP(6), B(5) => B_EXP(5), B(4) => B_EXP(4), 
                           B(3) => B_EXP(3), B(2) => B_EXP(2), B(1) => B_EXP(1)
                           , B(0) => B_EXP(0), CI => n1, SUM(7) => 
                           mw_I4sum_7_port, SUM(6) => EXP_in(6), SUM(5) => 
                           EXP_in(5), SUM(4) => EXP_in(4), SUM(3) => EXP_in(3),
                           SUM(2) => EXP_in(2), SUM(1) => EXP_in(1), SUM(0) => 
                           EXP_in(0), CO => n_1402, clk => clk);
   MY_CLK_r_REG1497_S1 : DFF_X1 port map( D => B_SIG(13), CK => clk, Q => n3800
                           , QN => n_1403);
   MY_CLK_r_REG1477_S1 : DFF_X1 port map( D => B_SIG(22), CK => clk, Q => n3804
                           , QN => n4679);
   MY_CLK_r_REG1502_S1 : DFF_X1 port map( D => B_SIG(11), CK => clk, Q => n3827
                           , QN => n_1404);
   MY_CLK_r_REG1040_S2 : DFF_X1 port map( D => mult_143_n5396, CK => clk, Q => 
                           n3701, QN => n_1405);
   MY_CLK_r_REG1215_S2 : DFF_X1 port map( D => n3022, CK => clk, Q => n3611, QN
                           => n_1406);
   MY_CLK_r_REG1368_S1 : DFF_X1 port map( D => mult_143_n4837, CK => clk, Q => 
                           n3553, QN => n_1407);
   MY_CLK_r_REG1475_S1 : DFF_X1 port map( D => B_SIG(22), CK => clk, Q => n3789
                           , QN => n_1408);
   MY_CLK_r_REG1450_S1 : DFF_X1 port map( D => mult_143_n3228, CK => clk, Q => 
                           n3536, QN => n_1409);
   MY_CLK_r_REG1441_S1 : DFF_X1 port map( D => n1738, CK => clk, Q => n3637, QN
                           => n_1410);
   MY_CLK_r_REG1232_S2 : DFF_X1 port map( D => mult_143_n5722, CK => clk, Q => 
                           n3708, QN => n_1411);
   MY_CLK_r_REG1213_S2 : DFF_X1 port map( D => n1558, CK => clk, Q => n3650, QN
                           => n_1412);
   MY_CLK_r_REG1184_S2 : DFF_X1 port map( D => n3016, CK => clk, Q => n3599, QN
                           => n_1413);
   MY_CLK_r_REG1181_S2 : DFF_X1 port map( D => n1684, CK => clk, Q => n3733, QN
                           => n_1414);
   MY_CLK_r_REG1041_S2 : DFF_X1 port map( D => n1697, CK => clk, Q => n3742, QN
                           => n_1415);
   MY_CLK_r_REG1482_S1 : DFF_X1 port map( D => B_SIG(19), CK => clk, Q => n3786
                           , QN => n4727);
   MY_CLK_r_REG1324_S1 : DFF_X1 port map( D => mult_143_n84, CK => clk, Q => 
                           n3540, QN => n4739);
   MY_CLK_r_REG1246_S1 : DFF_X1 port map( D => mult_143_n4891, CK => clk, Q => 
                           n3643, QN => n4631);
   MY_CLK_r_REG1247_S1 : DFF_X1 port map( D => mult_143_n96, CK => clk, Q => 
                           n3531, QN => n4622);
   MY_CLK_r_REG1478_S1 : DFF_X1 port map( D => B_SIG(21), CK => clk, Q => n3788
                           , QN => n4743);
   MY_CLK_r_REG1426_S1 : DFF_X1 port map( D => n1782, CK => clk, Q => n3803, QN
                           => n4657);
   U478 : BUF_X2 port map( A => n3790, Z => n4766);
   MY_CLK_r_REG1210_S3 : DFF_X1 port map( D => mult_143_n2755, CK => clk, Q => 
                           n3770, QN => n4612);
   U9 : CLKBUF_X1 port map( A => n3767, Z => n4665);
   U10 : CLKBUF_X1 port map( A => n1594, Z => n3120);
   U13 : CLKBUF_X1 port map( A => mult_143_n5389, Z => n4685);
   U18 : AOI222_X2 port map( A1 => mult_143_n5562, A2 => mult_143_n6402, B1 => 
                           mult_143_n5562, B2 => mult_143_n5564, C1 => 
                           mult_143_n6402, C2 => mult_143_n5564, ZN => 
                           mult_143_n5570);
   U136 : AOI222_X1 port map( A1 => n2755, A2 => n2606, B1 => n2755, B2 => 
                           mult_143_n4490, C1 => n2606, C2 => mult_143_n4490, 
                           ZN => mult_143_n5741);
   U305 : NAND2_X1 port map( A1 => mult_143_n2702, A2 => mult_143_n1719, ZN => 
                           n4980);
   U356 : XOR2_X1 port map( A => mult_143_n4984, B => mult_143_n4985, Z => 
                           n4981);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage1 is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         A_EXP : out std_logic_vector (7 downto 0);  A_SIG : out 
         std_logic_vector (31 downto 0);  B_EXP : out std_logic_vector (7 
         downto 0);  B_SIG : out std_logic_vector (31 downto 0);  
         SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : out 
         std_logic);

end FPmul_stage1;

architecture SYN_struct of FPmul_stage1 is

   component UnpackFP_1
      port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector
            (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, 
            isNaN, isINF, isZ, isDN : out std_logic);
   end component;
   
   component UnpackFP_0
      port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector
            (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, 
            isNaN, isINF, isZ, isDN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal A_isINF, A_isNaN, A_isZ, B_isINF, B_isNaN, B_isZ, A_SIGN, B_SIGN, n1,
      n2, n3, n4, n5, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449 : std_logic;

begin
   
   U11 : XOR2_X1 port map( A => B_SIGN, B => A_SIGN, Z => SIGN_out_stage1);
   U8 : NOR2_X1 port map( A1 => A_isNaN, A2 => B_isNaN, ZN => n3);
   U4 : OAI21_X1 port map( B1 => B_isZ, B2 => A_isZ, A => n3, ZN => n2);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => isZ_tab_stage1);
   U10 : NOR2_X1 port map( A1 => A_isINF, A2 => B_isINF, ZN => n5);
   U9 : AOI221_X1 port map( B1 => B_isZ, B2 => A_isINF, C1 => A_isZ, C2 => 
                           B_isINF, A => n5, ZN => isINF_stage1);
   U6 : AOI22_X1 port map( A1 => A_isINF, A2 => B_isZ, B1 => B_isINF, B2 => 
                           A_isZ, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n3, B2 => n1, A => n4, ZN => isNaN_stage1);
   U7 : OR2_X1 port map( A1 => A_isINF, A2 => B_isINF, ZN => n1);
   I0 : UnpackFP_0 port map( FP(31) => FP_A(31), FP(30) => FP_A(30), FP(29) => 
                           FP_A(29), FP(28) => FP_A(28), FP(27) => FP_A(27), 
                           FP(26) => FP_A(26), FP(25) => FP_A(25), FP(24) => 
                           FP_A(24), FP(23) => FP_A(23), FP(22) => FP_A(22), 
                           FP(21) => FP_A(21), FP(20) => FP_A(20), FP(19) => 
                           FP_A(19), FP(18) => FP_A(18), FP(17) => FP_A(17), 
                           FP(16) => FP_A(16), FP(15) => FP_A(15), FP(14) => 
                           FP_A(14), FP(13) => FP_A(13), FP(12) => FP_A(12), 
                           FP(11) => FP_A(11), FP(10) => FP_A(10), FP(9) => 
                           FP_A(9), FP(8) => FP_A(8), FP(7) => FP_A(7), FP(6) 
                           => FP_A(6), FP(5) => FP_A(5), FP(4) => FP_A(4), 
                           FP(3) => FP_A(3), FP(2) => FP_A(2), FP(1) => FP_A(1)
                           , FP(0) => FP_A(0), SIG(31) => n_1432, SIG(30) => 
                           n_1433, SIG(29) => n_1434, SIG(28) => n_1435, 
                           SIG(27) => n_1436, SIG(26) => n_1437, SIG(25) => 
                           n_1438, SIG(24) => n_1439, SIG(23) => A_SIG(23), 
                           SIG(22) => A_SIG(22), SIG(21) => A_SIG(21), SIG(20) 
                           => A_SIG(20), SIG(19) => A_SIG(19), SIG(18) => 
                           A_SIG(18), SIG(17) => A_SIG(17), SIG(16) => 
                           A_SIG(16), SIG(15) => A_SIG(15), SIG(14) => 
                           A_SIG(14), SIG(13) => A_SIG(13), SIG(12) => 
                           A_SIG(12), SIG(11) => A_SIG(11), SIG(10) => 
                           A_SIG(10), SIG(9) => A_SIG(9), SIG(8) => A_SIG(8), 
                           SIG(7) => A_SIG(7), SIG(6) => A_SIG(6), SIG(5) => 
                           A_SIG(5), SIG(4) => A_SIG(4), SIG(3) => A_SIG(3), 
                           SIG(2) => A_SIG(2), SIG(1) => A_SIG(1), SIG(0) => 
                           A_SIG(0), EXP(7) => A_EXP(7), EXP(6) => A_EXP(6), 
                           EXP(5) => A_EXP(5), EXP(4) => A_EXP(4), EXP(3) => 
                           A_EXP(3), EXP(2) => A_EXP(2), EXP(1) => A_EXP(1), 
                           EXP(0) => A_EXP(0), SIGN => A_SIGN, isNaN => A_isNaN
                           , isINF => A_isINF, isZ => A_isZ, isDN => n_1440);
   I1 : UnpackFP_1 port map( FP(31) => FP_B(31), FP(30) => FP_B(30), FP(29) => 
                           FP_B(29), FP(28) => FP_B(28), FP(27) => FP_B(27), 
                           FP(26) => FP_B(26), FP(25) => FP_B(25), FP(24) => 
                           FP_B(24), FP(23) => FP_B(23), FP(22) => FP_B(22), 
                           FP(21) => FP_B(21), FP(20) => FP_B(20), FP(19) => 
                           FP_B(19), FP(18) => FP_B(18), FP(17) => FP_B(17), 
                           FP(16) => FP_B(16), FP(15) => FP_B(15), FP(14) => 
                           FP_B(14), FP(13) => FP_B(13), FP(12) => FP_B(12), 
                           FP(11) => FP_B(11), FP(10) => FP_B(10), FP(9) => 
                           FP_B(9), FP(8) => FP_B(8), FP(7) => FP_B(7), FP(6) 
                           => FP_B(6), FP(5) => FP_B(5), FP(4) => FP_B(4), 
                           FP(3) => FP_B(3), FP(2) => FP_B(2), FP(1) => FP_B(1)
                           , FP(0) => FP_B(0), SIG(31) => n_1441, SIG(30) => 
                           n_1442, SIG(29) => n_1443, SIG(28) => n_1444, 
                           SIG(27) => n_1445, SIG(26) => n_1446, SIG(25) => 
                           n_1447, SIG(24) => n_1448, SIG(23) => B_SIG(23), 
                           SIG(22) => B_SIG(22), SIG(21) => B_SIG(21), SIG(20) 
                           => B_SIG(20), SIG(19) => B_SIG(19), SIG(18) => 
                           B_SIG(18), SIG(17) => B_SIG(17), SIG(16) => 
                           B_SIG(16), SIG(15) => B_SIG(15), SIG(14) => 
                           B_SIG(14), SIG(13) => B_SIG(13), SIG(12) => 
                           B_SIG(12), SIG(11) => B_SIG(11), SIG(10) => 
                           B_SIG(10), SIG(9) => B_SIG(9), SIG(8) => B_SIG(8), 
                           SIG(7) => B_SIG(7), SIG(6) => B_SIG(6), SIG(5) => 
                           B_SIG(5), SIG(4) => B_SIG(4), SIG(3) => B_SIG(3), 
                           SIG(2) => B_SIG(2), SIG(1) => B_SIG(1), SIG(0) => 
                           B_SIG(0), EXP(7) => B_EXP(7), EXP(6) => B_EXP(6), 
                           EXP(5) => B_EXP(5), EXP(4) => B_EXP(4), EXP(3) => 
                           B_EXP(3), EXP(2) => B_EXP(2), EXP(1) => B_EXP(1), 
                           EXP(0) => B_EXP(0), SIGN => B_SIGN, isNaN => B_isNaN
                           , isINF => B_isINF, isZ => B_isZ, isDN => n_1449);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         FP_Z : out std_logic_vector (31 downto 0));

end FPmul;

architecture SYN_pipeline of FPmul is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FPmul_stage4
      port( EXP_neg : in std_logic;  EXP_out_round : in std_logic_vector (7 
            downto 0);  EXP_pos, SIGN_out : in std_logic;  SIG_out_round : in 
            std_logic_vector (27 downto 0);  clk, isINF_tab, isNaN, isZ_tab : 
            in std_logic;  FP_Z : out std_logic_vector (31 downto 0));
   end component;
   
   component FPmul_stage3
      port( EXP_in : in std_logic_vector (7 downto 0);  EXP_neg_stage2, 
            EXP_pos_stage2, SIGN_out_stage2 : in std_logic;  SIG_in : in 
            std_logic_vector (27 downto 0);  clk, isINF_stage2, isNaN_stage2, 
            isZ_tab_stage2 : in std_logic;  EXP_neg : out std_logic;  
            EXP_out_round : out std_logic_vector (7 downto 0);  EXP_pos, 
            SIGN_out : out std_logic;  SIG_out_round : out std_logic_vector (27
            downto 0);  isINF_tab, isNaN, isZ_tab : out std_logic);
   end component;
   
   component FPmul_stage2
      port( A_EXP : in std_logic_vector (7 downto 0);  A_SIG : in 
            std_logic_vector (31 downto 0);  B_EXP : in std_logic_vector (7 
            downto 0);  B_SIG : in std_logic_vector (31 downto 0);  
            SIGN_out_stage1, clk, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : 
            in std_logic;  EXP_in : out std_logic_vector (7 downto 0);  
            EXP_neg_stage2, EXP_pos_stage2, SIGN_out_stage2 : out std_logic;  
            SIG_in : out std_logic_vector (27 downto 0);  isINF_stage2, 
            isNaN_stage2, isZ_tab_stage2 : out std_logic);
   end component;
   
   component FPmul_stage1
      port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic
            ;  A_EXP : out std_logic_vector (7 downto 0);  A_SIG : out 
            std_logic_vector (31 downto 0);  B_EXP : out std_logic_vector (7 
            downto 0);  B_SIG : out std_logic_vector (31 downto 0);  
            SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : out 
            std_logic);
   end component;
   
   signal A_EXP_7_port, A_EXP_6_port, A_EXP_5_port, A_EXP_4_port, A_EXP_3_port,
      A_EXP_2_port, A_EXP_1_port, A_EXP_0_port, A_SIG_23_port, A_SIG_22_port, 
      A_SIG_21_port, A_SIG_20_port, A_SIG_19_port, A_SIG_18_port, A_SIG_17_port
      , A_SIG_16_port, A_SIG_15_port, A_SIG_14_port, A_SIG_13_port, 
      A_SIG_12_port, A_SIG_11_port, A_SIG_10_port, A_SIG_9_port, A_SIG_8_port, 
      A_SIG_7_port, A_SIG_6_port, A_SIG_5_port, A_SIG_4_port, A_SIG_3_port, 
      A_SIG_2_port, A_SIG_1_port, A_SIG_0_port, B_EXP_7_port, B_EXP_6_port, 
      B_EXP_5_port, B_EXP_4_port, B_EXP_3_port, B_EXP_2_port, B_EXP_1_port, 
      B_EXP_0_port, B_SIG_22_port, B_SIG_21_port, B_SIG_20_port, B_SIG_19_port,
      B_SIG_18_port, B_SIG_17_port, B_SIG_16_port, B_SIG_15_port, B_SIG_14_port
      , B_SIG_13_port, B_SIG_12_port, B_SIG_11_port, B_SIG_10_port, 
      B_SIG_9_port, B_SIG_8_port, B_SIG_7_port, B_SIG_6_port, B_SIG_5_port, 
      B_SIG_4_port, B_SIG_3_port, B_SIG_2_port, B_SIG_1_port, B_SIG_0_port, 
      SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1, 
      EXP_in_7_port, EXP_in_6_port, EXP_in_5_port, EXP_in_4_port, EXP_in_3_port
      , EXP_in_2_port, EXP_in_1_port, EXP_in_0_port, EXP_neg_stage2, 
      EXP_pos_stage2, SIGN_out_stage2, SIG_in_27_port, SIG_in_26_port, 
      SIG_in_25_port, SIG_in_24_port, SIG_in_23_port, SIG_in_22_port, 
      SIG_in_21_port, SIG_in_20_port, SIG_in_19_port, SIG_in_18_port, 
      SIG_in_17_port, SIG_in_16_port, SIG_in_15_port, SIG_in_14_port, 
      SIG_in_13_port, SIG_in_12_port, SIG_in_11_port, SIG_in_10_port, 
      SIG_in_9_port, SIG_in_8_port, SIG_in_7_port, SIG_in_6_port, SIG_in_5_port
      , SIG_in_4_port, SIG_in_3_port, SIG_in_2_port, isINF_stage2, isNaN_stage2
      , isZ_tab_stage2, EXP_neg, EXP_out_round_7_port, EXP_out_round_6_port, 
      EXP_out_round_5_port, EXP_out_round_4_port, EXP_out_round_3_port, 
      EXP_out_round_2_port, EXP_out_round_1_port, EXP_out_round_0_port, EXP_pos
      , SIGN_out, SIG_out_round_26_port, SIG_out_round_25_port, 
      SIG_out_round_24_port, SIG_out_round_23_port, SIG_out_round_22_port, 
      SIG_out_round_21_port, SIG_out_round_20_port, SIG_out_round_19_port, 
      SIG_out_round_18_port, SIG_out_round_17_port, SIG_out_round_16_port, 
      SIG_out_round_15_port, SIG_out_round_14_port, SIG_out_round_13_port, 
      SIG_out_round_12_port, SIG_out_round_11_port, SIG_out_round_10_port, 
      SIG_out_round_9_port, SIG_out_round_8_port, SIG_out_round_7_port, 
      SIG_out_round_6_port, SIG_out_round_5_port, SIG_out_round_4_port, 
      SIG_out_round_3_port, isINF_tab, isNaN, isZ_tab, n1, n4, n5, n6, n7, n11,
      n12, n24, n22, n23, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, 
      n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, 
      n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473 : 
      std_logic;

begin
   
   n1 <= '0';
   n4 <= '0';
   n5 <= '0';
   n6 <= '0';
   n7 <= '0';
   I1 : FPmul_stage1 port map( FP_A(31) => FP_A(31), FP_A(30) => FP_A(30), 
                           FP_A(29) => FP_A(29), FP_A(28) => FP_A(28), FP_A(27)
                           => FP_A(27), FP_A(26) => FP_A(26), FP_A(25) => 
                           FP_A(25), FP_A(24) => FP_A(24), FP_A(23) => FP_A(23)
                           , FP_A(22) => FP_A(22), FP_A(21) => FP_A(21), 
                           FP_A(20) => FP_A(20), FP_A(19) => FP_A(19), FP_A(18)
                           => FP_A(18), FP_A(17) => FP_A(17), FP_A(16) => 
                           FP_A(16), FP_A(15) => FP_A(15), FP_A(14) => FP_A(14)
                           , FP_A(13) => FP_A(13), FP_A(12) => FP_A(12), 
                           FP_A(11) => FP_A(11), FP_A(10) => FP_A(10), FP_A(9) 
                           => FP_A(9), FP_A(8) => FP_A(8), FP_A(7) => FP_A(7), 
                           FP_A(6) => FP_A(6), FP_A(5) => FP_A(5), FP_A(4) => 
                           FP_A(4), FP_A(3) => FP_A(3), FP_A(2) => FP_A(2), 
                           FP_A(1) => FP_A(1), FP_A(0) => FP_A(0), FP_B(31) => 
                           FP_B(31), FP_B(30) => FP_B(30), FP_B(29) => FP_B(29)
                           , FP_B(28) => FP_B(28), FP_B(27) => FP_B(27), 
                           FP_B(26) => FP_B(26), FP_B(25) => FP_B(25), FP_B(24)
                           => FP_B(24), FP_B(23) => FP_B(23), FP_B(22) => 
                           FP_B(22), FP_B(21) => FP_B(21), FP_B(20) => FP_B(20)
                           , FP_B(19) => FP_B(19), FP_B(18) => FP_B(18), 
                           FP_B(17) => FP_B(17), FP_B(16) => FP_B(16), FP_B(15)
                           => FP_B(15), FP_B(14) => FP_B(14), FP_B(13) => 
                           FP_B(13), FP_B(12) => FP_B(12), FP_B(11) => FP_B(11)
                           , FP_B(10) => FP_B(10), FP_B(9) => FP_B(9), FP_B(8) 
                           => FP_B(8), FP_B(7) => FP_B(7), FP_B(6) => FP_B(6), 
                           FP_B(5) => FP_B(5), FP_B(4) => FP_B(4), FP_B(3) => 
                           FP_B(3), FP_B(2) => FP_B(2), FP_B(1) => FP_B(1), 
                           FP_B(0) => FP_B(0), clk => clk, A_EXP(7) => 
                           A_EXP_7_port, A_EXP(6) => A_EXP_6_port, A_EXP(5) => 
                           A_EXP_5_port, A_EXP(4) => A_EXP_4_port, A_EXP(3) => 
                           A_EXP_3_port, A_EXP(2) => A_EXP_2_port, A_EXP(1) => 
                           A_EXP_1_port, A_EXP(0) => A_EXP_0_port, A_SIG(31) =>
                           n_1450, A_SIG(30) => n_1451, A_SIG(29) => n_1452, 
                           A_SIG(28) => n_1453, A_SIG(27) => n_1454, A_SIG(26) 
                           => n_1455, A_SIG(25) => n_1456, A_SIG(24) => n_1457,
                           A_SIG(23) => A_SIG_23_port, A_SIG(22) => 
                           A_SIG_22_port, A_SIG(21) => A_SIG_21_port, A_SIG(20)
                           => A_SIG_20_port, A_SIG(19) => A_SIG_19_port, 
                           A_SIG(18) => A_SIG_18_port, A_SIG(17) => 
                           A_SIG_17_port, A_SIG(16) => A_SIG_16_port, A_SIG(15)
                           => A_SIG_15_port, A_SIG(14) => A_SIG_14_port, 
                           A_SIG(13) => A_SIG_13_port, A_SIG(12) => 
                           A_SIG_12_port, A_SIG(11) => A_SIG_11_port, A_SIG(10)
                           => A_SIG_10_port, A_SIG(9) => A_SIG_9_port, A_SIG(8)
                           => A_SIG_8_port, A_SIG(7) => A_SIG_7_port, A_SIG(6) 
                           => A_SIG_6_port, A_SIG(5) => A_SIG_5_port, A_SIG(4) 
                           => A_SIG_4_port, A_SIG(3) => A_SIG_3_port, A_SIG(2) 
                           => A_SIG_2_port, A_SIG(1) => A_SIG_1_port, A_SIG(0) 
                           => A_SIG_0_port, B_EXP(7) => B_EXP_7_port, B_EXP(6) 
                           => B_EXP_6_port, B_EXP(5) => B_EXP_5_port, B_EXP(4) 
                           => B_EXP_4_port, B_EXP(3) => B_EXP_3_port, B_EXP(2) 
                           => B_EXP_2_port, B_EXP(1) => B_EXP_1_port, B_EXP(0) 
                           => B_EXP_0_port, B_SIG(31) => n_1458, B_SIG(30) => 
                           n_1459, B_SIG(29) => n_1460, B_SIG(28) => n_1461, 
                           B_SIG(27) => n_1462, B_SIG(26) => n_1463, B_SIG(25) 
                           => n_1464, B_SIG(24) => n_1465, B_SIG(23) => n12, 
                           B_SIG(22) => B_SIG_22_port, B_SIG(21) => 
                           B_SIG_21_port, B_SIG(20) => B_SIG_20_port, B_SIG(19)
                           => B_SIG_19_port, B_SIG(18) => B_SIG_18_port, 
                           B_SIG(17) => B_SIG_17_port, B_SIG(16) => 
                           B_SIG_16_port, B_SIG(15) => B_SIG_15_port, B_SIG(14)
                           => B_SIG_14_port, B_SIG(13) => B_SIG_13_port, 
                           B_SIG(12) => B_SIG_12_port, B_SIG(11) => 
                           B_SIG_11_port, B_SIG(10) => B_SIG_10_port, B_SIG(9) 
                           => B_SIG_9_port, B_SIG(8) => B_SIG_8_port, B_SIG(7) 
                           => B_SIG_7_port, B_SIG(6) => B_SIG_6_port, B_SIG(5) 
                           => B_SIG_5_port, B_SIG(4) => B_SIG_4_port, B_SIG(3) 
                           => B_SIG_3_port, B_SIG(2) => B_SIG_2_port, B_SIG(1) 
                           => B_SIG_1_port, B_SIG(0) => B_SIG_0_port, 
                           SIGN_out_stage1 => SIGN_out_stage1, isINF_stage1 => 
                           isINF_stage1, isNaN_stage1 => isNaN_stage1, 
                           isZ_tab_stage1 => isZ_tab_stage1);
   I2 : FPmul_stage2 port map( A_EXP(7) => A_EXP_7_port, A_EXP(6) => 
                           A_EXP_6_port, A_EXP(5) => A_EXP_5_port, A_EXP(4) => 
                           A_EXP_4_port, A_EXP(3) => A_EXP_3_port, A_EXP(2) => 
                           A_EXP_2_port, A_EXP(1) => A_EXP_1_port, A_EXP(0) => 
                           A_EXP_0_port, A_SIG(31) => n1, A_SIG(30) => n1, 
                           A_SIG(29) => n1, A_SIG(28) => n1, A_SIG(27) => n1, 
                           A_SIG(26) => n1, A_SIG(25) => n1, A_SIG(24) => n1, 
                           A_SIG(23) => A_SIG_23_port, A_SIG(22) => 
                           A_SIG_22_port, A_SIG(21) => A_SIG_21_port, A_SIG(20)
                           => A_SIG_20_port, A_SIG(19) => A_SIG_19_port, 
                           A_SIG(18) => A_SIG_18_port, A_SIG(17) => 
                           A_SIG_17_port, A_SIG(16) => A_SIG_16_port, A_SIG(15)
                           => A_SIG_15_port, A_SIG(14) => A_SIG_14_port, 
                           A_SIG(13) => A_SIG_13_port, A_SIG(12) => 
                           A_SIG_12_port, A_SIG(11) => A_SIG_11_port, A_SIG(10)
                           => A_SIG_10_port, A_SIG(9) => A_SIG_9_port, A_SIG(8)
                           => A_SIG_8_port, A_SIG(7) => A_SIG_7_port, A_SIG(6) 
                           => A_SIG_6_port, A_SIG(5) => A_SIG_5_port, A_SIG(4) 
                           => A_SIG_4_port, A_SIG(3) => A_SIG_3_port, A_SIG(2) 
                           => A_SIG_2_port, A_SIG(1) => A_SIG_1_port, A_SIG(0) 
                           => A_SIG_0_port, B_EXP(7) => B_EXP_7_port, B_EXP(6) 
                           => B_EXP_6_port, B_EXP(5) => B_EXP_5_port, B_EXP(4) 
                           => B_EXP_4_port, B_EXP(3) => B_EXP_3_port, B_EXP(2) 
                           => B_EXP_2_port, B_EXP(1) => B_EXP_1_port, B_EXP(0) 
                           => B_EXP_0_port, B_SIG(31) => n1, B_SIG(30) => n1, 
                           B_SIG(29) => n1, B_SIG(28) => n1, B_SIG(27) => n1, 
                           B_SIG(26) => n1, B_SIG(25) => n1, B_SIG(24) => n1, 
                           B_SIG(23) => n12, B_SIG(22) => B_SIG_22_port, 
                           B_SIG(21) => B_SIG_21_port, B_SIG(20) => 
                           B_SIG_20_port, B_SIG(19) => B_SIG_19_port, B_SIG(18)
                           => B_SIG_18_port, B_SIG(17) => B_SIG_17_port, 
                           B_SIG(16) => B_SIG_16_port, B_SIG(15) => 
                           B_SIG_15_port, B_SIG(14) => B_SIG_14_port, B_SIG(13)
                           => B_SIG_13_port, B_SIG(12) => B_SIG_12_port, 
                           B_SIG(11) => B_SIG_11_port, B_SIG(10) => 
                           B_SIG_10_port, B_SIG(9) => B_SIG_9_port, B_SIG(8) =>
                           B_SIG_8_port, B_SIG(7) => B_SIG_7_port, B_SIG(6) => 
                           B_SIG_6_port, B_SIG(5) => B_SIG_5_port, B_SIG(4) => 
                           B_SIG_4_port, B_SIG(3) => B_SIG_3_port, B_SIG(2) => 
                           B_SIG_2_port, B_SIG(1) => B_SIG_1_port, B_SIG(0) => 
                           B_SIG_0_port, SIGN_out_stage1 => SIGN_out_stage1, 
                           clk => clk, isINF_stage1 => isINF_stage1, 
                           isNaN_stage1 => isNaN_stage1, isZ_tab_stage1 => 
                           isZ_tab_stage1, EXP_in(7) => EXP_in_7_port, 
                           EXP_in(6) => EXP_in_6_port, EXP_in(5) => 
                           EXP_in_5_port, EXP_in(4) => EXP_in_4_port, EXP_in(3)
                           => EXP_in_3_port, EXP_in(2) => EXP_in_2_port, 
                           EXP_in(1) => EXP_in_1_port, EXP_in(0) => 
                           EXP_in_0_port, EXP_neg_stage2 => EXP_neg_stage2, 
                           EXP_pos_stage2 => EXP_pos_stage2, SIGN_out_stage2 =>
                           SIGN_out_stage2, SIG_in(27) => SIG_in_27_port, 
                           SIG_in(26) => SIG_in_26_port, SIG_in(25) => 
                           SIG_in_25_port, SIG_in(24) => SIG_in_24_port, 
                           SIG_in(23) => SIG_in_23_port, SIG_in(22) => 
                           SIG_in_22_port, SIG_in(21) => SIG_in_21_port, 
                           SIG_in(20) => SIG_in_20_port, SIG_in(19) => 
                           SIG_in_19_port, SIG_in(18) => SIG_in_18_port, 
                           SIG_in(17) => SIG_in_17_port, SIG_in(16) => 
                           SIG_in_16_port, SIG_in(15) => SIG_in_15_port, 
                           SIG_in(14) => SIG_in_14_port, SIG_in(13) => 
                           SIG_in_13_port, SIG_in(12) => SIG_in_12_port, 
                           SIG_in(11) => SIG_in_11_port, SIG_in(10) => 
                           SIG_in_10_port, SIG_in(9) => SIG_in_9_port, 
                           SIG_in(8) => SIG_in_8_port, SIG_in(7) => 
                           SIG_in_7_port, SIG_in(6) => SIG_in_6_port, SIG_in(5)
                           => SIG_in_5_port, SIG_in(4) => SIG_in_4_port, 
                           SIG_in(3) => SIG_in_3_port, SIG_in(2) => 
                           SIG_in_2_port, SIG_in(1) => n_1466, SIG_in(0) => 
                           n_1467, isINF_stage2 => isINF_stage2, isNaN_stage2 
                           => isNaN_stage2, isZ_tab_stage2 => isZ_tab_stage2);
   I3 : FPmul_stage3 port map( EXP_in(7) => EXP_in_7_port, EXP_in(6) => 
                           EXP_in_6_port, EXP_in(5) => EXP_in_5_port, EXP_in(4)
                           => EXP_in_4_port, EXP_in(3) => EXP_in_3_port, 
                           EXP_in(2) => EXP_in_2_port, EXP_in(1) => 
                           EXP_in_1_port, EXP_in(0) => EXP_in_0_port, 
                           EXP_neg_stage2 => EXP_neg_stage2, EXP_pos_stage2 => 
                           EXP_pos_stage2, SIGN_out_stage2 => SIGN_out_stage2, 
                           SIG_in(27) => SIG_in_27_port, SIG_in(26) => 
                           SIG_in_26_port, SIG_in(25) => SIG_in_25_port, 
                           SIG_in(24) => SIG_in_24_port, SIG_in(23) => 
                           SIG_in_23_port, SIG_in(22) => SIG_in_22_port, 
                           SIG_in(21) => SIG_in_21_port, SIG_in(20) => 
                           SIG_in_20_port, SIG_in(19) => SIG_in_19_port, 
                           SIG_in(18) => SIG_in_18_port, SIG_in(17) => 
                           SIG_in_17_port, SIG_in(16) => SIG_in_16_port, 
                           SIG_in(15) => SIG_in_15_port, SIG_in(14) => 
                           SIG_in_14_port, SIG_in(13) => SIG_in_13_port, 
                           SIG_in(12) => SIG_in_12_port, SIG_in(11) => 
                           SIG_in_11_port, SIG_in(10) => SIG_in_10_port, 
                           SIG_in(9) => SIG_in_9_port, SIG_in(8) => 
                           SIG_in_8_port, SIG_in(7) => SIG_in_7_port, SIG_in(6)
                           => SIG_in_6_port, SIG_in(5) => SIG_in_5_port, 
                           SIG_in(4) => SIG_in_4_port, SIG_in(3) => 
                           SIG_in_3_port, SIG_in(2) => SIG_in_2_port, SIG_in(1)
                           => n4, SIG_in(0) => n5, clk => clk, isINF_stage2 => 
                           isINF_stage2, isNaN_stage2 => isNaN_stage2, 
                           isZ_tab_stage2 => isZ_tab_stage2, EXP_neg => EXP_neg
                           , EXP_out_round(7) => EXP_out_round_7_port, 
                           EXP_out_round(6) => EXP_out_round_6_port, 
                           EXP_out_round(5) => EXP_out_round_5_port, 
                           EXP_out_round(4) => EXP_out_round_4_port, 
                           EXP_out_round(3) => EXP_out_round_3_port, 
                           EXP_out_round(2) => EXP_out_round_2_port, 
                           EXP_out_round(1) => EXP_out_round_1_port, 
                           EXP_out_round(0) => EXP_out_round_0_port, EXP_pos =>
                           EXP_pos, SIGN_out => SIGN_out, SIG_out_round(27) => 
                           n11, SIG_out_round(26) => SIG_out_round_26_port, 
                           SIG_out_round(25) => SIG_out_round_25_port, 
                           SIG_out_round(24) => SIG_out_round_24_port, 
                           SIG_out_round(23) => SIG_out_round_23_port, 
                           SIG_out_round(22) => SIG_out_round_22_port, 
                           SIG_out_round(21) => SIG_out_round_21_port, 
                           SIG_out_round(20) => SIG_out_round_20_port, 
                           SIG_out_round(19) => SIG_out_round_19_port, 
                           SIG_out_round(18) => SIG_out_round_18_port, 
                           SIG_out_round(17) => SIG_out_round_17_port, 
                           SIG_out_round(16) => SIG_out_round_16_port, 
                           SIG_out_round(15) => SIG_out_round_15_port, 
                           SIG_out_round(14) => SIG_out_round_14_port, 
                           SIG_out_round(13) => SIG_out_round_13_port, 
                           SIG_out_round(12) => SIG_out_round_12_port, 
                           SIG_out_round(11) => SIG_out_round_11_port, 
                           SIG_out_round(10) => SIG_out_round_10_port, 
                           SIG_out_round(9) => SIG_out_round_9_port, 
                           SIG_out_round(8) => SIG_out_round_8_port, 
                           SIG_out_round(7) => SIG_out_round_7_port, 
                           SIG_out_round(6) => SIG_out_round_6_port, 
                           SIG_out_round(5) => SIG_out_round_5_port, 
                           SIG_out_round(4) => SIG_out_round_4_port, 
                           SIG_out_round(3) => SIG_out_round_3_port, 
                           SIG_out_round(2) => n_1468, SIG_out_round(1) => 
                           n_1469, SIG_out_round(0) => n_1470, isINF_tab => 
                           isINF_tab, isNaN => isNaN, isZ_tab => isZ_tab);
   I4 : FPmul_stage4 port map( EXP_neg => EXP_neg, EXP_out_round(7) => 
                           EXP_out_round_7_port, EXP_out_round(6) => 
                           EXP_out_round_6_port, EXP_out_round(5) => 
                           EXP_out_round_5_port, EXP_out_round(4) => 
                           EXP_out_round_4_port, EXP_out_round(3) => 
                           EXP_out_round_3_port, EXP_out_round(2) => 
                           EXP_out_round_2_port, EXP_out_round(1) => 
                           EXP_out_round_1_port, EXP_out_round(0) => 
                           EXP_out_round_0_port, EXP_pos => EXP_pos, SIGN_out 
                           => SIGN_out, SIG_out_round(27) => n11, 
                           SIG_out_round(26) => SIG_out_round_26_port, 
                           SIG_out_round(25) => SIG_out_round_25_port, 
                           SIG_out_round(24) => SIG_out_round_24_port, 
                           SIG_out_round(23) => SIG_out_round_23_port, 
                           SIG_out_round(22) => SIG_out_round_22_port, 
                           SIG_out_round(21) => SIG_out_round_21_port, 
                           SIG_out_round(20) => SIG_out_round_20_port, 
                           SIG_out_round(19) => SIG_out_round_19_port, 
                           SIG_out_round(18) => SIG_out_round_18_port, 
                           SIG_out_round(17) => SIG_out_round_17_port, 
                           SIG_out_round(16) => SIG_out_round_16_port, 
                           SIG_out_round(15) => SIG_out_round_15_port, 
                           SIG_out_round(14) => SIG_out_round_14_port, 
                           SIG_out_round(13) => SIG_out_round_13_port, 
                           SIG_out_round(12) => SIG_out_round_12_port, 
                           SIG_out_round(11) => SIG_out_round_11_port, 
                           SIG_out_round(10) => SIG_out_round_10_port, 
                           SIG_out_round(9) => SIG_out_round_9_port, 
                           SIG_out_round(8) => SIG_out_round_8_port, 
                           SIG_out_round(7) => SIG_out_round_7_port, 
                           SIG_out_round(6) => SIG_out_round_6_port, 
                           SIG_out_round(5) => SIG_out_round_5_port, 
                           SIG_out_round(4) => SIG_out_round_4_port, 
                           SIG_out_round(3) => SIG_out_round_3_port, 
                           SIG_out_round(2) => n1, SIG_out_round(1) => n6, 
                           SIG_out_round(0) => n7, clk => clk, isINF_tab => 
                           isINF_tab, isNaN => isNaN, isZ_tab => isZ_tab, 
                           FP_Z(31) => n24, FP_Z(30) => FP_Z(30), FP_Z(29) => 
                           FP_Z(29), FP_Z(28) => FP_Z(28), FP_Z(27) => FP_Z(27)
                           , FP_Z(26) => FP_Z(26), FP_Z(25) => FP_Z(25), 
                           FP_Z(24) => FP_Z(24), FP_Z(23) => FP_Z(23), FP_Z(22)
                           => FP_Z(22), FP_Z(21) => FP_Z(21), FP_Z(20) => 
                           FP_Z(20), FP_Z(19) => FP_Z(19), FP_Z(18) => FP_Z(18)
                           , FP_Z(17) => FP_Z(17), FP_Z(16) => FP_Z(16), 
                           FP_Z(15) => FP_Z(15), FP_Z(14) => FP_Z(14), FP_Z(13)
                           => FP_Z(13), FP_Z(12) => FP_Z(12), FP_Z(11) => 
                           FP_Z(11), FP_Z(10) => FP_Z(10), FP_Z(9) => FP_Z(9), 
                           FP_Z(8) => FP_Z(8), FP_Z(7) => FP_Z(7), FP_Z(6) => 
                           FP_Z(6), FP_Z(5) => FP_Z(5), FP_Z(4) => FP_Z(4), 
                           FP_Z(3) => FP_Z(3), FP_Z(2) => FP_Z(2), FP_Z(1) => 
                           FP_Z(1), FP_Z(0) => FP_Z(0));
   MY_CLK_r_REG1023_S5 : DFF_X1 port map( D => n22, CK => clk, Q => FP_Z(31), 
                           QN => n_1471);
   MY_CLK_r_REG1022_S4 : DFF_X1 port map( D => n23, CK => clk, Q => n22, QN => 
                           n_1472);
   MY_CLK_r_REG1021_S3 : DFF_X1 port map( D => n24, CK => clk, Q => n23, QN => 
                           n_1473);

end SYN_pipeline;
