package my_pkg is

	constant n_levels : 6;

end my_pkg;
