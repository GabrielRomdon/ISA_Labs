
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_FPmul is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_FPmul;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         FP_Z : out std_logic_vector (31 downto 0));

end FPmul;

architecture SYN_pipeline of FPmul is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFRS_X1
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SDFF_X2
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal A_EXP_7_port, A_EXP_6_port, A_EXP_5_port, A_EXP_4_port, A_EXP_3_port,
      A_EXP_2_port, A_EXP_1_port, A_EXP_0_port, A_SIG_23_port, A_SIG_16_port, 
      A_SIG_10_port, A_SIG_8_port, B_EXP_7_port, B_EXP_6_port, B_EXP_5_port, 
      B_EXP_4_port, B_EXP_3_port, B_EXP_2_port, B_EXP_1_port, B_EXP_0_port, 
      B_SIG_9_port, B_SIG_8_port, SIGN_out_stage1, isINF_stage1, isNaN_stage1, 
      isZ_tab_stage1, EXP_in_7_port, EXP_in_5_port, EXP_in_3_port, 
      EXP_in_2_port, EXP_neg_stage2, EXP_pos_stage2, SIGN_out_stage2, 
      SIG_in_27_port, SIG_in_26_port, SIG_in_11_port, SIG_in_4_port, 
      SIG_in_3_port, isINF_stage2, isNaN_stage2, isZ_tab_stage2, EXP_neg, 
      EXP_out_round_7_port, EXP_out_round_5_port, EXP_out_round_4_port, 
      EXP_out_round_3_port, EXP_out_round_2_port, EXP_out_round_1_port, 
      SIG_out_round_26_port, SIG_out_round_25_port, isINF_tab, I1_isZ_tab_int, 
      I1_isNaN_int, I1_isINF_int, I1_SIGN_out_int, I2_dtemp_23_port, 
      I2_dtemp_26_port, I2_dtemp_27_port, I2_dtemp_28_port, I2_dtemp_30_port, 
      I2_dtemp_31_port, I2_dtemp_33_port, I2_dtemp_34_port, I2_dtemp_37_port, 
      I2_dtemp_38_port, I2_dtemp_39_port, I2_dtemp_40_port, I2_dtemp_41_port, 
      I2_dtemp_42_port, I2_dtemp_43_port, I2_dtemp_44_port, I2_mw_I4sum_0_port,
      I2_mw_I4sum_1_port, I2_mw_I4sum_2_port, I2_mw_I4sum_3_port, 
      I2_mw_I4sum_4_port, I2_mw_I4sum_5_port, I2_mw_I4sum_6_port, I2_N0, 
      I2_SIGN_out_stage2_tmp, I2_isZ_tab_stage2_tmp, I2_isNaN_stage2_tmp, 
      I2_isINF_stage2_tmp, I2_EXP_neg_stage2_tmp, I2_EXP_pos_int, 
      I2_EXP_pos_stage2_tmp, I2_EXP_in_tmp_0_port, I2_EXP_in_tmp_1_port, 
      I2_EXP_in_tmp_2_port, I2_EXP_in_tmp_3_port, I2_EXP_in_tmp_5_port, 
      I2_EXP_in_tmp_6_port, I2_EXP_in_tmp_7_port, I2_SIG_in_int_2_port, 
      I2_SIG_in_int_3_port, I2_SIG_in_int_4_port, I2_SIG_in_int_5_port, 
      I2_SIG_in_int_6_port, I2_SIG_in_int_7_port, I2_SIG_in_int_8_port, 
      I2_SIG_in_int_9_port, I2_SIG_in_int_10_port, I2_SIG_in_int_11_port, 
      I2_SIG_in_int_12_port, I2_SIG_in_int_13_port, I2_SIG_in_int_14_port, 
      I2_SIG_in_int_15_port, I2_SIG_in_int_16_port, I2_SIG_in_int_17_port, 
      I2_SIG_in_int_18_port, I2_SIG_in_int_19_port, I2_SIG_in_int_20_port, 
      I2_SIG_in_int_21_port, I2_SIG_in_int_22_port, I2_SIG_in_int_23_port, 
      I2_SIG_in_int_24_port, I2_SIG_in_int_25_port, I2_SIG_in_int_26_port, 
      I2_SIG_in_int_27_port, I3_SIG_out_3_port, I3_SIG_out_4_port, 
      I3_SIG_out_5_port, I3_SIG_out_6_port, I3_SIG_out_7_port, 
      I3_SIG_out_8_port, I3_SIG_out_9_port, I3_SIG_out_10_port, 
      I3_SIG_out_11_port, I3_SIG_out_12_port, I3_SIG_out_13_port, 
      I3_SIG_out_14_port, I3_SIG_out_15_port, I3_SIG_out_16_port, 
      I3_SIG_out_17_port, I3_SIG_out_18_port, I3_SIG_out_19_port, 
      I3_SIG_out_20_port, I3_SIG_out_21_port, I3_SIG_out_22_port, 
      I3_SIG_out_23_port, I3_SIG_out_24_port, I3_SIG_out_25_port, 
      I3_SIG_out_27_port, I3_EXP_out_0_port, I3_EXP_out_1_port, 
      I3_EXP_out_2_port, I3_EXP_out_3_port, I3_EXP_out_4_port, 
      I3_EXP_out_5_port, I3_EXP_out_6_port, I3_EXP_out_7_port, I4_FP_0_port, 
      I4_FP_1_port, I4_FP_2_port, I4_FP_3_port, I4_FP_4_port, I4_FP_5_port, 
      I4_FP_6_port, I4_FP_7_port, I4_FP_8_port, I4_FP_9_port, I4_FP_10_port, 
      I4_FP_11_port, I4_FP_12_port, I4_FP_13_port, I4_FP_14_port, I4_FP_15_port
      , I4_FP_16_port, I4_FP_17_port, I4_FP_18_port, I4_FP_19_port, 
      I4_FP_20_port, I4_FP_21_port, I4_FP_22_port, I4_FP_23_port, I4_FP_24_port
      , I4_FP_25_port, I4_FP_26_port, I4_FP_27_port, I4_FP_28_port, 
      I4_FP_29_port, I4_FP_30_port, I4_FP_31_port, I1_I0_N13, I1_I1_N13, 
      mult_x_19_n4, n164, n200, n204, n205, n356, n357, n358, n359, n360, n362,
      n363, n364, n365, n366, n367, n369, n370, n371, n372, n373, n374, n376, 
      n377, n379, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n2555, n2556, n2557, n2558, n2559, n2560, 
      n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, 
      n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2579, n2582, n2583, 
      n2584, n2587, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, 
      n2597, n2598, n2599, n2600, n2601, n2602, n2604, n2605, n2606, n2608, 
      n2611, n2613, n2638, intadd_33_A_1_port, intadd_33_A_0_port, 
      intadd_33_B_2_port, intadd_33_B_1_port, intadd_33_B_0_port, intadd_33_CI,
      intadd_33_SUM_2_port, intadd_33_SUM_1_port, intadd_33_SUM_0_port, 
      intadd_33_n3, intadd_33_n2, intadd_33_n1, intadd_2_CI, intadd_2_n6, 
      intadd_2_n5, intadd_2_n4, intadd_2_n3, intadd_2_n2, intadd_2_n1, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4356, n4357, n4358, 
      n4359, n4360, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, 
      n4370, n4371, n4372, n4373, n4374, n4375, n4377, n4378, n4379, n4380, 
      n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4389, n4390, n4391, 
      n4392, n4393, n4395, n4396, n4397, n4398, n4399, n4401, n4402, n4403, 
      n4405, n4406, n4407, n4408, n4409, n4411, n4412, n4413, n4414, n4415, 
      n4416, n4417, n4418, n4420, n4421, n4422, n4423, n4424, n4425, n4426, 
      n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, 
      n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4447, n4448, 
      n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
      n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4467, n4468, n4469, 
      n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, 
      n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4489, n4490, 
      n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, 
      n4501, n4503, n4504, n4506, n4507, n4508, n4509, n4510, n4511, n4512, 
      n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4522, n4523, n4524, 
      n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, 
      n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, 
      n4545, n4546, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, 
      n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, 
      n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, 
      n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, 
      n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, 
      n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, 
      n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, 
      n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, 
      n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, 
      n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, 
      n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, 
      n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, 
      n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, 
      n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, 
      n4686, n4687, n4688, n4689, n4690, n4691, n4693, n4694, n4695, n4696, 
      n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, 
      n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, 
      n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, 
      n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4736, n4737, 
      n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, 
      n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
      n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, 
      n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, 
      n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, 
      n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, 
      n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, 
      n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, 
      n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, 
      n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, 
      n4838, n4839, n4840, n4841, n4843, n4844, n4845, n4846, n4847, n4848, 
      n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, 
      n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, 
      n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, 
      n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, 
      n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, 
      n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, 
      n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, 
      n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, 
      n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, 
      n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, 
      n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, 
      n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, 
      n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, 
      n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, 
      n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4997, n4998, n4999, 
      n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, 
      n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, 
      n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, 
      n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, 
      n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, 
      n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, 
      n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, 
      n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, 
      n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, 
      n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, 
      n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, 
      n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, 
      n5121, n5122, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, 
      n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, 
      n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, 
      n5152, n5153, n5154, n5155, n5156, n5158, n5159, n5160, n5161, n5162, 
      n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, 
      n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, 
      n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, 
      n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, 
      n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, 
      n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, 
      n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, 
      n5233, n5234, n5235, n5237, n5238, n5239, n5240, n5241, n5242, n5243, 
      n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, 
      n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, 
      n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, 
      n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, 
      n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, 
      n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, 
      n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, 
      n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, 
      n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, 
      n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, 
      n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, 
      n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, 
      n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, 
      n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, 
      n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, 
      n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, 
      n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5436, 
      n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, 
      n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, 
      n5457, n5458, n5459, n5460, n5461, n5463, n5464, n5465, n5466, n5467, 
      n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, 
      n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, 
      n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, 
      n5498, n5499, n5500, n5501, n5502, n5504, n5505, n5506, n5507, n5508, 
      n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, 
      n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, 
      n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, 
      n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, 
      n5549, n5550, n5551, n5553, n5554, n5555, n5557, n5558, n5559, n5560, 
      n5561, n5562, n5563, n5564, n5565, n5566, n5568, n5569, n5570, n5571, 
      n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, 
      n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, 
      n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, 
      n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, 
      n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, 
      n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, 
      n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, 
      n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, 
      n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, 
      n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, 
      n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, 
      n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, 
      n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, 
      n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, 
      n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, 
      n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, 
      n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, 
      n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, 
      n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, 
      n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, 
      n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, 
      n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, 
      n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, 
      n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, 
      n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, 
      n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, 
      n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
      n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, 
      n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
      n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, 
      n5883, n5884, n5885, n5886, n5887, n5889, n5890, n5891, n5892, n5893, 
      n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, 
      n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, 
      n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, 
      n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, 
      n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, 
      n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, 
      n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, 
      n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, 
      n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, 
      n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, 
      n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, 
      n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, 
      n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, 
      n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, 
      n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, 
      n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, 
      n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, 
      n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, 
      n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, 
      n6085, n6086, n6087, n6089, n6090, n6091, n6092, n6093, n6094, n6095, 
      n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, 
      n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6116, 
      n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, 
      n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, 
      n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, 
      n6169, n6170, n6171, n6172, n6174, n6175, n6176, n6177, n6178, n6179, 
      n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, 
      n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, 
      n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, 
      n6210, n6211, n6212, n6213, n6214, n6215, n6217, n6218, n6219, n6220, 
      n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, 
      n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6242, 
      n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, 
      n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, 
      n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, 
      n6273, n6274, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, 
      n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, 
      n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, 
      n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, 
      n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, 
      n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, 
      n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, 
      n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, 
      n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, 
      n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, 
      n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, 
      n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, 
      n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, 
      n6405, n6406, n6407, n6408, n6409, n6411, n6412, n6413, n6414, n6415, 
      n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, 
      n6427, n6428, n6429, n6430, n6431, n6433, n6434, n6435, n6436, n6437, 
      n6438, n6439, n6440, n6441, n6442, n6443, n6445, n6446, n6447, n6448, 
      n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, 
      n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6469, 
      n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, 
      n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, 
      n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, 
      n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6509, n6510, 
      n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6521, n6522, 
      n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, 
      n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, 
      n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, 
      n6553, n6554, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, 
      n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, 
      n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, 
      n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, 
      n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6605, 
      n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, 
      n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, 
      n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, 
      n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6645, n6646, 
      n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, 
      n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, 
      n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, 
      n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6686, n6687, 
      n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6698, 
      n6699, n6700, n6701, n6702, n6703, n6705, n6706, n6707, n6708, n6709, 
      n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, 
      n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, 
      n6730, n6731, n6732, n6733, n6734, n6736, n6737, n6738, n6739, n6740, 
      n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, 
      n6751, n6752, n6753, n6754, n6756, n6757, n6758, n6759, n6760, n6761, 
      n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, 
      n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, 
      n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6791, n6792, 
      n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, 
      n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, 
      n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, 
      n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, 
      n6834, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, 
      n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, 
      n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, 
      n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
      n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
      n6886, n6887, n6888, n6889, n6891, n6892, n6893, n6894, n6895, n6896, 
      n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, 
      n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, 
      n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, 
      n6927, n6928, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, 
      n6938, n6939, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, 
      n6949, n6950, n6951, n6953, n6954, n6955, n6956, n6957, n6958, n6959, 
      n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, 
      n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, 
      n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, 
      n6990, n6991, n6992, n6994, n6995, n6996, n6997, n6998, n6999, n7000, 
      n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, 
      n7011, n7012, n7013, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
      n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7030, n7031, n7032, 
      n7033, n7034, n7035, n7036, n7038, n7039, n7040, n7041, n7042, n7043, 
      n7044, n7045, n7046, n7047, n7048, n7049, n7051, n7052, n7053, n7054, 
      n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, 
      n7065, n7066, n7067, n7068, n7069, n7070, n7073, n7074, n7075, n7076, 
      n7077, n7078, n7079, n7080, n7081, n7082, n7084, n7085, n7086, n7087, 
      n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, 
      n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, 
      n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7117, n7118, 
      n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, 
      n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, 
      n7139, n7140, n7141, n7144, n7145, n7146, n7147, n7148, n7149, n7150, 
      n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, 
      n7161, n7162, n7163, n7164, n7165, n7167, n7168, n7169, n7170, n7171, 
      n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, 
      n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, 
      n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, 
      n7202, n7203, n7204, n7205, n7206, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, 
      n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, 
      n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, 
      n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, 
      n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, 
      n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, 
      n7355, n7356, n7357, n7358, n7359, n7360, n7362, n7363, n7364, n7365, 
      n7366, n7367, n7368, n7370, n7371, n7372, n7373, n7374, n7375, n7376, 
      n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, 
      n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, 
      n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, 
      n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, 
      n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, 
      n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, 
      n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, 
      n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, 
      n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, 
      n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, 
      n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, 
      n7488, n7489, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, 
      n7499, n7500, n7501, n7503, n7504, n7505, n7506, n7508, n7509, n7510, 
      n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, 
      n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, 
      n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, 
      n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, 
      n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, 
      n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, 
      n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7582, 
      n7583, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7623, n7624, 
      n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, 
      n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, 
      n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, 
      n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, 
      n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, 
      n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, 
      n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, 
      n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, 
      n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, 
      n7715, n7716, n7717, n7718, n7719, n7721, n7722, n7723, n7724, n7725, 
      n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, 
      n7737, n7738, n7739, n7740, n7742, n7743, n7744, n7745, n7746, n7747, 
      n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, 
      n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, 
      n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, 
      n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, 
      n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, 
      n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, 
      n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, 
      n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, 
      n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, 
      n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, 
      n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, 
      n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, 
      n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, 
      n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, 
      n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, 
      n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, 
      n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, 
      n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, 
      n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, 
      n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, 
      n7948, n7949, n7951, n7952, n7953, n7955, n7956, n7957, n7958, n7959, 
      n7960, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, 
      n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, 
      n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7991, 
      n7992, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, 
      n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, 
      n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, 
      n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, 
      n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, 
      n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, 
      n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, 
      n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, 
      n8073, n8074, n8075, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
      n8094, n8095, n8096, n8098, n8099, n8100, n8101, n8102, n8103, n8104, 
      n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, 
      n8115, n8116, n8117, n8118, n8119, n8121, n8122, n8123, n8124, n8125, 
      n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8134, n8135, n8136, 
      n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, 
      n8147, n8148, n8149, n8150, n8152, n8154, n8155, n8156, n8157, n8158, 
      n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, 
      n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, 
      n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, 
      n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8198, n8199, 
      n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, 
      n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, 
      n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, 
      n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, 
      n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, 
      n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, 
      n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, 
      n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, 
      n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, 
      n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, 
      n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, 
      n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8323, n8324, 
      n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, 
      n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, 
      n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, 
      n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, 
      n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, 
      n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, 
      n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, 
      n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8403, n8404, n8405, 
      n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, 
      n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, 
      n8426, n8428, n8429, n8430, n8431, n8434, n8436, n8438, n8441, n8443, 
      n8444, n8445, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, 
      n8456, n8458, n8459, n8461, n8462, n8464, n8465, n8466, n8467, n8468, 
      n8469, n8470, n8471, n8472, n8473, n8474, n8476, n8478, n8479, n8480, 
      n8481, n8484, n8485, n8487, n8488, n8489, n8490, n8492, n8495, n8496, 
      n8497, n8498, n8500, n8501, n8502, n8503, n8504, n8506, n8510, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8520, n8522, n8526, n8527, n8528, 
      n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, 
      n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, 
      n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, 
      n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, 
      n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, 
      n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, 
      n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, 
      n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, 
      n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, 
      n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, 
      n8629, n8630, n8631, n8632, n_1000, n_1001, n_1002, n_1003, n_1004, 
      n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, 
      n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, 
      n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, 
      n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, 
      n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, 
      n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, 
      n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, 
      n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, 
      n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, 
      n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, 
      n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, 
      n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, 
      n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, 
      n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, 
      n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, 
      n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, 
      n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, 
      n_1158 : std_logic;

begin
   
   I1_B_SIG_reg_5_inst : DFF_X1 port map( D => FP_B(5), CK => clk, Q => n8401, 
                           QN => n376);
   I1_B_EXP_reg_0_inst : DFF_X1 port map( D => FP_B(23), CK => clk, Q => 
                           B_EXP_0_port, QN => n8382);
   I1_B_EXP_reg_1_inst : DFF_X1 port map( D => FP_B(24), CK => clk, Q => 
                           B_EXP_1_port, QN => n_1000);
   I1_B_EXP_reg_2_inst : DFF_X1 port map( D => FP_B(25), CK => clk, Q => 
                           B_EXP_2_port, QN => n_1001);
   I1_B_EXP_reg_4_inst : DFF_X1 port map( D => FP_B(27), CK => clk, Q => 
                           B_EXP_4_port, QN => n_1002);
   I1_B_EXP_reg_5_inst : DFF_X1 port map( D => FP_B(28), CK => clk, Q => 
                           B_EXP_5_port, QN => n_1003);
   I1_B_EXP_reg_6_inst : DFF_X1 port map( D => FP_B(29), CK => clk, Q => 
                           B_EXP_6_port, QN => n_1004);
   I1_B_EXP_reg_7_inst : DFF_X1 port map( D => FP_B(30), CK => clk, Q => 
                           B_EXP_7_port, QN => n_1005);
   I1_isNaN_stage1_reg : DFF_X1 port map( D => I1_isNaN_int, CK => clk, Q => 
                           isNaN_stage1, QN => n_1006);
   I1_isINF_stage1_reg : DFF_X1 port map( D => I1_isINF_int, CK => clk, Q => 
                           isINF_stage1, QN => n_1007);
   I1_A_SIG_reg_2_inst : DFF_X1 port map( D => FP_A(2), CK => clk, Q => n8370, 
                           QN => n366);
   I1_A_SIG_reg_3_inst : DFF_X1 port map( D => FP_A(3), CK => clk, Q => n8356, 
                           QN => n392);
   I1_A_SIG_reg_4_inst : DFF_X1 port map( D => FP_A(4), CK => clk, Q => n8363, 
                           QN => n367);
   I1_A_SIG_reg_6_inst : DFF_X1 port map( D => FP_A(6), CK => clk, Q => n8335, 
                           QN => n164);
   I1_A_SIG_reg_8_inst : DFF_X1 port map( D => FP_A(8), CK => clk, Q => 
                           A_SIG_8_port, QN => n8368);
   I1_A_SIG_reg_10_inst : DFF_X1 port map( D => FP_A(10), CK => clk, Q => 
                           A_SIG_10_port, QN => n8366);
   I1_A_SIG_reg_12_inst : DFF_X1 port map( D => FP_A(12), CK => clk, Q => n8360
                           , QN => n369);
   I1_A_SIG_reg_14_inst : DFF_X1 port map( D => FP_A(14), CK => clk, Q => n8361
                           , QN => n358);
   I1_A_SIG_reg_16_inst : DFF_X1 port map( D => FP_A(16), CK => clk, Q => 
                           A_SIG_16_port, QN => n8357);
   I1_A_SIG_reg_18_inst : DFF_X1 port map( D => FP_A(18), CK => clk, Q => n8359
                           , QN => n365);
   I1_A_SIG_reg_20_inst : DFF_X1 port map( D => FP_A(20), CK => clk, Q => n8400
                           , QN => n370);
   I1_A_SIG_reg_22_inst : DFF_X1 port map( D => FP_A(22), CK => clk, Q => n8364
                           , QN => n200);
   I1_A_SIG_reg_23_inst : DFF_X1 port map( D => I1_I0_N13, CK => clk, Q => 
                           A_SIG_23_port, QN => n8398);
   I1_A_EXP_reg_0_inst : DFF_X1 port map( D => FP_A(23), CK => clk, Q => 
                           A_EXP_0_port, QN => n8344);
   I1_A_EXP_reg_1_inst : DFF_X1 port map( D => FP_A(24), CK => clk, Q => 
                           A_EXP_1_port, QN => n_1008);
   I1_A_EXP_reg_2_inst : DFF_X1 port map( D => FP_A(25), CK => clk, Q => 
                           A_EXP_2_port, QN => n_1009);
   I1_A_EXP_reg_3_inst : DFF_X1 port map( D => FP_A(26), CK => clk, Q => 
                           A_EXP_3_port, QN => n_1010);
   I1_A_EXP_reg_4_inst : DFF_X1 port map( D => FP_A(27), CK => clk, Q => 
                           A_EXP_4_port, QN => n_1011);
   I1_A_EXP_reg_5_inst : DFF_X1 port map( D => FP_A(28), CK => clk, Q => 
                           A_EXP_5_port, QN => n_1012);
   I1_A_EXP_reg_6_inst : DFF_X1 port map( D => FP_A(29), CK => clk, Q => 
                           A_EXP_6_port, QN => n_1013);
   I1_A_EXP_reg_7_inst : DFF_X1 port map( D => FP_A(30), CK => clk, Q => 
                           A_EXP_7_port, QN => n_1014);
   I1_SIGN_out_stage1_reg : DFF_X1 port map( D => I1_SIGN_out_int, CK => clk, Q
                           => SIGN_out_stage1, QN => n_1015);
   I2_prod_tmp_reg_22_inst : DFF_X1 port map( D => n8407, CK => clk, Q => 
                           I2_SIG_in_int_2_port, QN => n_1016);
   I2_prod_tmp_reg_27_inst : DFF_X1 port map( D => I2_dtemp_27_port, CK => clk,
                           Q => I2_SIG_in_int_7_port, QN => n_1017);
   I2_prod_tmp_reg_29_inst : DFF_X1 port map( D => n8406, CK => clk, Q => 
                           I2_SIG_in_int_9_port, QN => n_1018);
   I2_prod_tmp_reg_33_inst : DFF_X1 port map( D => I2_dtemp_33_port, CK => clk,
                           Q => I2_SIG_in_int_13_port, QN => n_1019);
   I2_prod_tmp_reg_34_inst : DFF_X1 port map( D => I2_dtemp_34_port, CK => clk,
                           Q => I2_SIG_in_int_14_port, QN => n_1020);
   I2_prod_tmp_reg_35_inst : DFF_X1 port map( D => n8410, CK => clk, Q => 
                           I2_SIG_in_int_15_port, QN => n_1021);
   I2_prod_tmp_reg_37_inst : DFF_X1 port map( D => I2_dtemp_37_port, CK => clk,
                           Q => I2_SIG_in_int_17_port, QN => n_1022);
   I2_prod_tmp_reg_43_inst : DFF_X1 port map( D => I2_dtemp_43_port, CK => clk,
                           Q => I2_SIG_in_int_23_port, QN => n_1023);
   I2_SIGN_out_stage2_tmp_reg : DFF_X1 port map( D => SIGN_out_stage1, CK => 
                           clk, Q => I2_SIGN_out_stage2_tmp, QN => n_1024);
   I2_SIGN_out_stage2_reg : DFF_X1 port map( D => I2_SIGN_out_stage2_tmp, CK =>
                           clk, Q => SIGN_out_stage2, QN => n_1025);
   I2_isZ_tab_stage2_tmp_reg : DFF_X1 port map( D => isZ_tab_stage1, CK => clk,
                           Q => I2_isZ_tab_stage2_tmp, QN => n_1026);
   I2_isZ_tab_stage2_reg : DFF_X1 port map( D => I2_isZ_tab_stage2_tmp, CK => 
                           clk, Q => isZ_tab_stage2, QN => n_1027);
   I2_isNaN_stage2_tmp_reg : DFF_X1 port map( D => isNaN_stage1, CK => clk, Q 
                           => I2_isNaN_stage2_tmp, QN => n_1028);
   I2_isNaN_stage2_reg : DFF_X1 port map( D => I2_isNaN_stage2_tmp, CK => clk, 
                           Q => isNaN_stage2, QN => n_1029);
   I2_isINF_stage2_tmp_reg : DFF_X1 port map( D => isINF_stage1, CK => clk, Q 
                           => I2_isINF_stage2_tmp, QN => n_1030);
   I2_isINF_stage2_reg : DFF_X1 port map( D => I2_isINF_stage2_tmp, CK => clk, 
                           Q => isINF_stage2, QN => n_1031);
   I2_EXP_neg_stage2_tmp_reg : DFF_X1 port map( D => I2_N0, CK => clk, Q => 
                           I2_EXP_neg_stage2_tmp, QN => n_1032);
   I2_EXP_neg_stage2_reg : DFF_X1 port map( D => I2_EXP_neg_stage2_tmp, CK => 
                           clk, Q => EXP_neg_stage2, QN => n_1033);
   I2_EXP_pos_stage2_tmp_reg : DFF_X1 port map( D => I2_EXP_pos_int, CK => clk,
                           Q => I2_EXP_pos_stage2_tmp, QN => n_1034);
   I2_EXP_pos_stage2_reg : DFF_X1 port map( D => I2_EXP_pos_stage2_tmp, CK => 
                           clk, Q => EXP_pos_stage2, QN => n_1035);
   I2_SIG_in_reg_3_inst : DFF_X1 port map( D => I2_SIG_in_int_3_port, CK => clk
                           , Q => SIG_in_3_port, QN => n_1036);
   I2_SIG_in_reg_4_inst : DFF_X1 port map( D => I2_SIG_in_int_4_port, CK => clk
                           , Q => SIG_in_4_port, QN => n8373);
   I2_SIG_in_reg_5_inst : DFF_X1 port map( D => I2_SIG_in_int_5_port, CK => clk
                           , Q => n_1037, QN => n8341);
   I2_SIG_in_reg_6_inst : DFF_X1 port map( D => I2_SIG_in_int_6_port, CK => clk
                           , Q => n_1038, QN => n2608);
   I2_SIG_in_reg_7_inst : DFF_X1 port map( D => I2_SIG_in_int_7_port, CK => clk
                           , Q => n_1039, QN => n8365);
   I2_SIG_in_reg_8_inst : DFF_X1 port map( D => I2_SIG_in_int_8_port, CK => clk
                           , Q => n_1040, QN => n2606);
   I2_SIG_in_reg_9_inst : DFF_X1 port map( D => I2_SIG_in_int_9_port, CK => clk
                           , Q => n8381, QN => n2605);
   I2_SIG_in_reg_10_inst : DFF_X1 port map( D => I2_SIG_in_int_10_port, CK => 
                           clk, Q => n8371, QN => n2604);
   I2_SIG_in_reg_11_inst : DFF_X1 port map( D => I2_SIG_in_int_11_port, CK => 
                           clk, Q => SIG_in_11_port, QN => n8374);
   I2_SIG_in_reg_12_inst : DFF_X1 port map( D => I2_SIG_in_int_12_port, CK => 
                           clk, Q => n_1041, QN => n2602);
   I2_SIG_in_reg_13_inst : DFF_X1 port map( D => I2_SIG_in_int_13_port, CK => 
                           clk, Q => n8345, QN => n2601);
   I2_SIG_in_reg_14_inst : DFF_X1 port map( D => I2_SIG_in_int_14_port, CK => 
                           clk, Q => n8387, QN => n2600);
   I2_SIG_in_reg_15_inst : DFF_X1 port map( D => I2_SIG_in_int_15_port, CK => 
                           clk, Q => n8346, QN => n2599);
   I2_SIG_in_reg_16_inst : DFF_X1 port map( D => I2_SIG_in_int_16_port, CK => 
                           clk, Q => n8388, QN => n2598);
   I2_SIG_in_reg_17_inst : DFF_X1 port map( D => I2_SIG_in_int_17_port, CK => 
                           clk, Q => n_1042, QN => n2597);
   I2_SIG_in_reg_18_inst : DFF_X1 port map( D => I2_SIG_in_int_18_port, CK => 
                           clk, Q => n_1043, QN => n2596);
   I2_SIG_in_reg_22_inst : DFF_X1 port map( D => I2_SIG_in_int_22_port, CK => 
                           clk, Q => n_1044, QN => n2592);
   I2_SIG_in_reg_23_inst : DFF_X1 port map( D => I2_SIG_in_int_23_port, CK => 
                           clk, Q => n8347, QN => n2591);
   I2_SIG_in_reg_24_inst : DFF_X1 port map( D => I2_SIG_in_int_24_port, CK => 
                           clk, Q => n8389, QN => n2590);
   I2_SIG_in_reg_25_inst : DFF_X1 port map( D => I2_SIG_in_int_25_port, CK => 
                           clk, Q => n8380, QN => n2589);
   I2_EXP_in_tmp_reg_0_inst : DFF_X1 port map( D => I2_mw_I4sum_0_port, CK => 
                           clk, Q => I2_EXP_in_tmp_0_port, QN => n_1045);
   I2_EXP_in_tmp_reg_1_inst : DFF_X1 port map( D => I2_mw_I4sum_1_port, CK => 
                           clk, Q => I2_EXP_in_tmp_1_port, QN => n_1046);
   I2_EXP_in_reg_1_inst : DFF_X1 port map( D => I2_EXP_in_tmp_1_port, CK => clk
                           , Q => n_1047, QN => n2577);
   I2_EXP_in_tmp_reg_2_inst : DFF_X1 port map( D => I2_mw_I4sum_2_port, CK => 
                           clk, Q => I2_EXP_in_tmp_2_port, QN => n_1048);
   I2_EXP_in_reg_2_inst : DFF_X1 port map( D => I2_EXP_in_tmp_2_port, CK => clk
                           , Q => EXP_in_2_port, QN => n_1049);
   I2_EXP_in_tmp_reg_3_inst : DFF_X1 port map( D => I2_mw_I4sum_3_port, CK => 
                           clk, Q => I2_EXP_in_tmp_3_port, QN => n_1050);
   I2_EXP_in_reg_3_inst : DFF_X1 port map( D => I2_EXP_in_tmp_3_port, CK => clk
                           , Q => EXP_in_3_port, QN => n8343);
   I2_EXP_in_tmp_reg_5_inst : DFF_X1 port map( D => I2_mw_I4sum_5_port, CK => 
                           clk, Q => I2_EXP_in_tmp_5_port, QN => n_1051);
   I2_EXP_in_reg_5_inst : DFF_X1 port map( D => I2_EXP_in_tmp_5_port, CK => clk
                           , Q => EXP_in_5_port, QN => n8384);
   I2_EXP_in_tmp_reg_6_inst : DFF_X1 port map( D => I2_mw_I4sum_6_port, CK => 
                           clk, Q => I2_EXP_in_tmp_6_port, QN => n_1052);
   I2_EXP_in_reg_6_inst : DFF_X1 port map( D => I2_EXP_in_tmp_6_port, CK => clk
                           , Q => n8376, QN => n_1053);
   I2_EXP_in_tmp_reg_7_inst : DFF_X1 port map( D => n374, CK => clk, Q => 
                           I2_EXP_in_tmp_7_port, QN => n_1054);
   I2_EXP_in_reg_7_inst : DFF_X1 port map( D => I2_EXP_in_tmp_7_port, CK => clk
                           , Q => EXP_in_7_port, QN => n_1055);
   I3_EXP_neg_reg : DFF_X1 port map( D => EXP_neg_stage2, CK => clk, Q => 
                           EXP_neg, QN => n_1056);
   I3_EXP_pos_reg : DFF_X1 port map( D => EXP_pos_stage2, CK => clk, Q => 
                           n_1057, QN => n2613);
   I3_SIGN_out_reg : DFF_X1 port map( D => SIGN_out_stage2, CK => clk, Q => 
                           I4_FP_31_port, QN => n_1058);
   I3_isZ_tab_reg : DFF_X1 port map( D => isZ_tab_stage2, CK => clk, Q => 
                           n_1059, QN => n2611);
   I3_isNaN_reg : DFF_X1 port map( D => isNaN_stage2, CK => clk, Q => n_1060, 
                           QN => n2567);
   I3_isINF_tab_reg : DFF_X1 port map( D => isINF_stage2, CK => clk, Q => 
                           isINF_tab, QN => n8385);
   I3_SIG_out_round_reg_3_inst : DFF_X1 port map( D => I3_SIG_out_3_port, CK =>
                           clk, Q => n_1061, QN => n2587);
   I3_SIG_out_round_reg_4_inst : DFF_X1 port map( D => I3_SIG_out_4_port, CK =>
                           clk, Q => n_1062, QN => n2565);
   I3_SIG_out_round_reg_5_inst : DFF_X1 port map( D => I3_SIG_out_5_port, CK =>
                           clk, Q => n_1063, QN => n2556);
   I3_SIG_out_round_reg_6_inst : DFF_X1 port map( D => I3_SIG_out_6_port, CK =>
                           clk, Q => n_1064, QN => n2568);
   I3_SIG_out_round_reg_7_inst : DFF_X1 port map( D => I3_SIG_out_7_port, CK =>
                           clk, Q => n_1065, QN => n2557);
   I3_SIG_out_round_reg_8_inst : DFF_X1 port map( D => I3_SIG_out_8_port, CK =>
                           clk, Q => n_1066, QN => n2569);
   I3_SIG_out_round_reg_9_inst : DFF_X1 port map( D => I3_SIG_out_9_port, CK =>
                           clk, Q => n_1067, QN => n2558);
   I3_SIG_out_round_reg_10_inst : DFF_X1 port map( D => I3_SIG_out_10_port, CK 
                           => clk, Q => n_1068, QN => n2570);
   I3_SIG_out_round_reg_11_inst : DFF_X1 port map( D => I3_SIG_out_11_port, CK 
                           => clk, Q => n_1069, QN => n2559);
   I3_SIG_out_round_reg_12_inst : DFF_X1 port map( D => I3_SIG_out_12_port, CK 
                           => clk, Q => n_1070, QN => n2571);
   I3_SIG_out_round_reg_13_inst : DFF_X1 port map( D => I3_SIG_out_13_port, CK 
                           => clk, Q => n_1071, QN => n2560);
   I3_SIG_out_round_reg_14_inst : DFF_X1 port map( D => I3_SIG_out_14_port, CK 
                           => clk, Q => n_1072, QN => n2572);
   I3_SIG_out_round_reg_15_inst : DFF_X1 port map( D => I3_SIG_out_15_port, CK 
                           => clk, Q => n_1073, QN => n2561);
   I3_SIG_out_round_reg_16_inst : DFF_X1 port map( D => I3_SIG_out_16_port, CK 
                           => clk, Q => n_1074, QN => n2573);
   I3_SIG_out_round_reg_17_inst : DFF_X1 port map( D => I3_SIG_out_17_port, CK 
                           => clk, Q => n_1075, QN => n2562);
   I3_SIG_out_round_reg_18_inst : DFF_X1 port map( D => I3_SIG_out_18_port, CK 
                           => clk, Q => n_1076, QN => n2574);
   I3_SIG_out_round_reg_19_inst : DFF_X1 port map( D => I3_SIG_out_19_port, CK 
                           => clk, Q => n_1077, QN => n2563);
   I3_SIG_out_round_reg_20_inst : DFF_X1 port map( D => I3_SIG_out_20_port, CK 
                           => clk, Q => n_1078, QN => n2575);
   I3_SIG_out_round_reg_21_inst : DFF_X1 port map( D => I3_SIG_out_21_port, CK 
                           => clk, Q => n_1079, QN => n2564);
   I3_SIG_out_round_reg_22_inst : DFF_X1 port map( D => I3_SIG_out_22_port, CK 
                           => clk, Q => n_1080, QN => n2576);
   I3_SIG_out_round_reg_23_inst : DFF_X1 port map( D => I3_SIG_out_23_port, CK 
                           => clk, Q => n_1081, QN => n2555);
   I3_SIG_out_round_reg_24_inst : DFF_X1 port map( D => I3_SIG_out_24_port, CK 
                           => clk, Q => n_1082, QN => n2566);
   I3_SIG_out_round_reg_25_inst : DFF_X1 port map( D => I3_SIG_out_25_port, CK 
                           => clk, Q => SIG_out_round_25_port, QN => n8342);
   I3_SIG_out_round_reg_27_inst : DFF_X1 port map( D => I3_SIG_out_27_port, CK 
                           => clk, Q => n8377, QN => n2582);
   I3_EXP_out_round_reg_0_inst : DFF_X1 port map( D => I3_EXP_out_0_port, CK =>
                           clk, Q => n_1083, QN => n2584);
   I3_EXP_out_round_reg_1_inst : DFF_X1 port map( D => I3_EXP_out_1_port, CK =>
                           clk, Q => EXP_out_round_1_port, QN => n_1084);
   I3_EXP_out_round_reg_2_inst : DFF_X1 port map( D => I3_EXP_out_2_port, CK =>
                           clk, Q => EXP_out_round_2_port, QN => n8390);
   I3_EXP_out_round_reg_3_inst : DFF_X1 port map( D => I3_EXP_out_3_port, CK =>
                           clk, Q => EXP_out_round_3_port, QN => n_1085);
   I3_EXP_out_round_reg_4_inst : DFF_X1 port map( D => I3_EXP_out_4_port, CK =>
                           clk, Q => EXP_out_round_4_port, QN => n_1086);
   I3_EXP_out_round_reg_5_inst : DFF_X1 port map( D => I3_EXP_out_5_port, CK =>
                           clk, Q => EXP_out_round_5_port, QN => n8379);
   I3_EXP_out_round_reg_6_inst : DFF_X1 port map( D => I3_EXP_out_6_port, CK =>
                           clk, Q => n8383, QN => n2579);
   I4_FP_Z_reg_0_inst : DFF_X1 port map( D => I4_FP_0_port, CK => clk, Q => 
                           FP_Z(0), QN => n_1087);
   I4_FP_Z_reg_1_inst : DFF_X1 port map( D => I4_FP_1_port, CK => clk, Q => 
                           FP_Z(1), QN => n_1088);
   I4_FP_Z_reg_2_inst : DFF_X1 port map( D => I4_FP_2_port, CK => clk, Q => 
                           FP_Z(2), QN => n_1089);
   I4_FP_Z_reg_3_inst : DFF_X1 port map( D => I4_FP_3_port, CK => clk, Q => 
                           FP_Z(3), QN => n_1090);
   I4_FP_Z_reg_4_inst : DFF_X1 port map( D => I4_FP_4_port, CK => clk, Q => 
                           FP_Z(4), QN => n_1091);
   I4_FP_Z_reg_5_inst : DFF_X1 port map( D => I4_FP_5_port, CK => clk, Q => 
                           FP_Z(5), QN => n_1092);
   I4_FP_Z_reg_6_inst : DFF_X1 port map( D => I4_FP_6_port, CK => clk, Q => 
                           FP_Z(6), QN => n_1093);
   I4_FP_Z_reg_7_inst : DFF_X1 port map( D => I4_FP_7_port, CK => clk, Q => 
                           FP_Z(7), QN => n_1094);
   I4_FP_Z_reg_8_inst : DFF_X1 port map( D => I4_FP_8_port, CK => clk, Q => 
                           FP_Z(8), QN => n_1095);
   I4_FP_Z_reg_9_inst : DFF_X1 port map( D => I4_FP_9_port, CK => clk, Q => 
                           FP_Z(9), QN => n_1096);
   I4_FP_Z_reg_10_inst : DFF_X1 port map( D => I4_FP_10_port, CK => clk, Q => 
                           FP_Z(10), QN => n_1097);
   I4_FP_Z_reg_11_inst : DFF_X1 port map( D => I4_FP_11_port, CK => clk, Q => 
                           FP_Z(11), QN => n_1098);
   I4_FP_Z_reg_12_inst : DFF_X1 port map( D => I4_FP_12_port, CK => clk, Q => 
                           FP_Z(12), QN => n_1099);
   I4_FP_Z_reg_13_inst : DFF_X1 port map( D => I4_FP_13_port, CK => clk, Q => 
                           FP_Z(13), QN => n_1100);
   I4_FP_Z_reg_14_inst : DFF_X1 port map( D => I4_FP_14_port, CK => clk, Q => 
                           FP_Z(14), QN => n_1101);
   I4_FP_Z_reg_15_inst : DFF_X1 port map( D => I4_FP_15_port, CK => clk, Q => 
                           FP_Z(15), QN => n_1102);
   I4_FP_Z_reg_16_inst : DFF_X1 port map( D => I4_FP_16_port, CK => clk, Q => 
                           FP_Z(16), QN => n_1103);
   I4_FP_Z_reg_17_inst : DFF_X1 port map( D => I4_FP_17_port, CK => clk, Q => 
                           FP_Z(17), QN => n_1104);
   I4_FP_Z_reg_18_inst : DFF_X1 port map( D => I4_FP_18_port, CK => clk, Q => 
                           FP_Z(18), QN => n_1105);
   I4_FP_Z_reg_19_inst : DFF_X1 port map( D => I4_FP_19_port, CK => clk, Q => 
                           FP_Z(19), QN => n_1106);
   I4_FP_Z_reg_20_inst : DFF_X1 port map( D => I4_FP_20_port, CK => clk, Q => 
                           FP_Z(20), QN => n_1107);
   I4_FP_Z_reg_21_inst : DFF_X1 port map( D => I4_FP_21_port, CK => clk, Q => 
                           FP_Z(21), QN => n_1108);
   I4_FP_Z_reg_22_inst : DFF_X1 port map( D => I4_FP_22_port, CK => clk, Q => 
                           FP_Z(22), QN => n_1109);
   I4_FP_Z_reg_23_inst : DFF_X1 port map( D => I4_FP_23_port, CK => clk, Q => 
                           FP_Z(23), QN => n_1110);
   I4_FP_Z_reg_24_inst : DFF_X1 port map( D => I4_FP_24_port, CK => clk, Q => 
                           FP_Z(24), QN => n_1111);
   I4_FP_Z_reg_25_inst : DFF_X1 port map( D => I4_FP_25_port, CK => clk, Q => 
                           FP_Z(25), QN => n_1112);
   I4_FP_Z_reg_26_inst : DFF_X1 port map( D => I4_FP_26_port, CK => clk, Q => 
                           FP_Z(26), QN => n_1113);
   I4_FP_Z_reg_27_inst : DFF_X1 port map( D => I4_FP_27_port, CK => clk, Q => 
                           FP_Z(27), QN => n_1114);
   I4_FP_Z_reg_28_inst : DFF_X1 port map( D => I4_FP_28_port, CK => clk, Q => 
                           FP_Z(28), QN => n_1115);
   I4_FP_Z_reg_29_inst : DFF_X1 port map( D => I4_FP_29_port, CK => clk, Q => 
                           FP_Z(29), QN => n_1116);
   I4_FP_Z_reg_30_inst : DFF_X1 port map( D => I4_FP_30_port, CK => clk, Q => 
                           FP_Z(30), QN => n_1117);
   I4_FP_Z_reg_31_inst : DFF_X1 port map( D => I4_FP_31_port, CK => clk, Q => 
                           FP_Z(31), QN => n_1118);
   I1_isZ_tab_stage1_reg : DFF_X1 port map( D => I1_isZ_tab_int, CK => clk, Q 
                           => isZ_tab_stage1, QN => n_1119);
   I1_A_SIG_reg_0_inst : DFF_X1 port map( D => FP_A(0), CK => clk, Q => n8358, 
                           QN => mult_x_19_n4);
   I1_B_SIG_reg_23_inst : DFF_X1 port map( D => I1_I1_N13, CK => clk, Q => 
                           n8336, QN => n364);
   I2_prod_tmp_reg_24_inst : DFF_X1 port map( D => n8414, CK => clk, Q => 
                           I2_SIG_in_int_4_port, QN => n_1120);
   I3_EXP_out_round_reg_7_inst : DFF_X1 port map( D => I3_EXP_out_7_port, CK =>
                           clk, Q => EXP_out_round_7_port, QN => n_1121);
   I2_prod_tmp_reg_46_inst : DFF_X1 port map( D => n8412, CK => clk, Q => 
                           I2_SIG_in_int_26_port, QN => n_1122);
   I2_prod_tmp_reg_42_inst : DFF_X1 port map( D => I2_dtemp_42_port, CK => clk,
                           Q => I2_SIG_in_int_22_port, QN => n_1123);
   I2_prod_tmp_reg_36_inst : DFF_X1 port map( D => n8409, CK => clk, Q => 
                           I2_SIG_in_int_16_port, QN => n_1124);
   I2_prod_tmp_reg_45_inst : DFF_X1 port map( D => n8411, CK => clk, Q => 
                           I2_SIG_in_int_25_port, QN => n_1125);
   I2_prod_tmp_reg_25_inst : DFF_X1 port map( D => n8413, CK => clk, Q => 
                           I2_SIG_in_int_5_port, QN => n_1126);
   I2_prod_tmp_reg_23_inst : DFF_X1 port map( D => I2_dtemp_23_port, CK => clk,
                           Q => I2_SIG_in_int_3_port, QN => n_1127);
   I1_B_SIG_reg_8_inst : DFF_X1 port map( D => FP_B(8), CK => clk, Q => 
                           B_SIG_8_port, QN => n8362);
   intadd_33_U4 : FA_X1 port map( A => intadd_33_A_0_port, B => 
                           intadd_33_B_0_port, CI => intadd_33_CI, CO => 
                           intadd_33_n3, S => intadd_33_SUM_0_port);
   intadd_33_U3 : FA_X1 port map( A => intadd_33_A_1_port, B => 
                           intadd_33_B_1_port, CI => intadd_33_n3, CO => 
                           intadd_33_n2, S => intadd_33_SUM_1_port);
   intadd_33_U2 : FA_X1 port map( A => n8408, B => intadd_33_B_2_port, CI => 
                           intadd_33_n2, CO => intadd_33_n1, S => 
                           intadd_33_SUM_2_port);
   intadd_2_U7 : FA_X1 port map( A => A_EXP_1_port, B => B_EXP_1_port, CI => 
                           intadd_2_CI, CO => intadd_2_n6, S => 
                           I2_mw_I4sum_1_port);
   intadd_2_U6 : FA_X1 port map( A => A_EXP_2_port, B => B_EXP_2_port, CI => 
                           intadd_2_n6, CO => intadd_2_n5, S => 
                           I2_mw_I4sum_2_port);
   intadd_2_U5 : FA_X1 port map( A => A_EXP_3_port, B => B_EXP_3_port, CI => 
                           intadd_2_n5, CO => intadd_2_n4, S => 
                           I2_mw_I4sum_3_port);
   intadd_2_U4 : FA_X1 port map( A => A_EXP_4_port, B => B_EXP_4_port, CI => 
                           intadd_2_n4, CO => intadd_2_n3, S => 
                           I2_mw_I4sum_4_port);
   intadd_2_U3 : FA_X1 port map( A => A_EXP_5_port, B => B_EXP_5_port, CI => 
                           intadd_2_n3, CO => intadd_2_n2, S => 
                           I2_mw_I4sum_5_port);
   intadd_2_U2 : FA_X1 port map( A => A_EXP_6_port, B => B_EXP_6_port, CI => 
                           intadd_2_n2, CO => intadd_2_n1, S => 
                           I2_mw_I4sum_6_port);
   I1_A_SIG_reg_21_inst : DFF_X1 port map( D => FP_A(21), CK => clk, Q => n8399
                           , QN => n387);
   I1_A_SIG_reg_1_inst : DFF_X1 port map( D => FP_A(1), CK => clk, Q => n8395, 
                           QN => n385);
   I1_A_SIG_reg_17_inst : DFF_X1 port map( D => FP_A(17), CK => clk, Q => n8353
                           , QN => n383);
   I1_A_SIG_reg_7_inst : DFF_X1 port map( D => FP_A(7), CK => clk, Q => n8355, 
                           QN => n389);
   I1_A_SIG_reg_9_inst : DFF_X1 port map( D => FP_A(9), CK => clk, Q => n8338, 
                           QN => n388);
   I1_A_SIG_reg_11_inst : DFF_X1 port map( D => FP_A(11), CK => clk, Q => n8340
                           , QN => n382);
   I1_A_SIG_reg_15_inst : DFF_X1 port map( D => FP_A(15), CK => clk, Q => n8369
                           , QN => n384);
   I1_A_SIG_reg_19_inst : DFF_X1 port map( D => FP_A(19), CK => clk, Q => n8339
                           , QN => n393);
   I1_B_SIG_reg_0_inst : DFF_X2 port map( D => FP_B(0), CK => clk, Q => n8354, 
                           QN => n2638);
   I1_B_SIG_reg_11_inst : DFF_X2 port map( D => FP_B(11), CK => clk, Q => n8392
                           , QN => n379);
   I1_B_SIG_reg_4_inst : DFF_X2 port map( D => FP_B(4), CK => clk, Q => n8350, 
                           QN => n8324);
   I1_B_SIG_reg_14_inst : DFF_X2 port map( D => FP_B(14), CK => clk, Q => n8394
                           , QN => n359);
   I1_B_SIG_reg_17_inst : DFF_X2 port map( D => FP_B(17), CK => clk, Q => n8330
                           , QN => n372);
   I1_B_SIG_reg_9_inst : DFF_X2 port map( D => FP_B(9), CK => clk, Q => 
                           B_SIG_9_port, QN => n8327);
   I1_B_SIG_reg_10_inst : DFF_X2 port map( D => FP_B(10), CK => clk, Q => n8351
                           , QN => n204);
   I2_SIG_in_reg_26_inst : DFF_X1 port map( D => I2_SIG_in_int_26_port, CK => 
                           clk, Q => SIG_in_26_port, QN => n8375);
   I2_EXP_in_reg_0_inst : DFF_X1 port map( D => I2_EXP_in_tmp_0_port, CK => clk
                           , Q => n8386, QN => n2583);
   I2_SIG_in_reg_21_inst : DFF_X1 port map( D => I2_SIG_in_int_21_port, CK => 
                           clk, Q => n_1128, QN => n2593);
   I2_SIG_in_reg_19_inst : DFF_X1 port map( D => I2_SIG_in_int_19_port, CK => 
                           clk, Q => n8391, QN => n2595);
   I1_A_SIG_reg_5_inst : DFF_X1 port map( D => FP_A(5), CK => clk, Q => n8397, 
                           QN => n391);
   I1_A_SIG_reg_13_inst : DFF_X1 port map( D => FP_A(13), CK => clk, Q => n8403
                           , QN => n394);
   I1_B_SIG_reg_22_inst : SDFF_X2 port map( D => n8317, SI => n8318, SE => 
                           FP_B(22), CK => clk, Q => n357, QN => n8331);
   I1_B_SIG_reg_21_inst : DFF_X1 port map( D => FP_B(21), CK => clk, Q => n8334
                           , QN => n205);
   I1_B_SIG_reg_1_inst : DFF_X1 port map( D => FP_B(1), CK => clk, Q => n8393, 
                           QN => n395);
   I1_B_SIG_reg_19_inst : DFF_X1 port map( D => FP_B(19), CK => clk, Q => n8325
                           , QN => n371);
   I1_B_SIG_reg_13_inst : DFF_X1 port map( D => FP_B(13), CK => clk, Q => n8326
                           , QN => n356);
   I1_B_SIG_reg_16_inst : DFF_X2 port map( D => FP_B(16), CK => clk, Q => n8337
                           , QN => n360);
   U1730 : XNOR2_X1 port map( A => n5735, B => n5734, ZN => n6073);
   U1732 : NAND2_X1 port map( A1 => n4350, A2 => n4349, ZN => n5252);
   U1734 : NAND2_X1 port map( A1 => n5173, A2 => n5172, ZN => n4349);
   U1735 : INV_X1 port map( A => n4750, ZN => n4659);
   U1738 : NAND3_X1 port map( A1 => n7972, A2 => n7971, A3 => n7974, ZN => 
                           n7980);
   U1742 : INV_X1 port map( A => n6121, ZN => n6118);
   U1744 : NAND2_X1 port map( A1 => n4347, A2 => n4531, ZN => n4522);
   U1747 : XNOR2_X1 port map( A => n5515, B => n5514, ZN => n5553);
   U1752 : XNOR2_X1 port map( A => n4348, B => n8150, ZN => I2_dtemp_34_port);
   U1753 : NAND3_X1 port map( A1 => n8184, A2 => n8480, A3 => n8192, ZN => 
                           n4348);
   U1754 : NAND2_X2 port map( A1 => n4892, A2 => n8358, ZN => n7946);
   U1756 : NAND2_X1 port map( A1 => n4657, A2 => n4656, ZN => n4750);
   U1762 : OAI21_X1 port map( B1 => n5173, B2 => n5172, A => n5171, ZN => n4350
                           );
   U1772 : NAND2_X1 port map( A1 => n6151, A2 => n4352, ZN => n6157);
   U1773 : NAND2_X1 port map( A1 => n6153, A2 => n6152, ZN => n4352);
   U1775 : NAND2_X1 port map( A1 => n7215, A2 => n8423, ZN => n4353);
   U1778 : NAND2_X1 port map( A1 => n7195, A2 => n4381, ZN => n4380);
   U1779 : NAND2_X1 port map( A1 => n7105, A2 => n7104, ZN => n7191);
   U1780 : INV_X1 port map( A => n7692, ZN => n5746);
   U1781 : NAND2_X1 port map( A1 => n5114, A2 => n5113, ZN => n4356);
   U1782 : XNOR2_X2 port map( A => n7184, B => n7265, ZN => n4443);
   U1783 : AND3_X1 port map( A1 => n4459, A2 => n8254, A3 => n8223, ZN => n4357
                           );
   U1784 : AND2_X1 port map( A1 => n7591, A2 => n7590, ZN => n4358);
   U1785 : AND3_X1 port map( A1 => n8252, A2 => n8601, A3 => n8223, ZN => n4359
                           );
   U1786 : NAND2_X1 port map( A1 => n8514, A2 => n8403, ZN => n4360);
   U1787 : NAND2_X1 port map( A1 => n4962, A2 => n8403, ZN => n7120);
   U1789 : AND4_X1 port map( A1 => n7480, A2 => n8585, A3 => n7636, A4 => n7601
                           , ZN => n4417);
   U1796 : INV_X1 port map( A => n4379, ZN => n8092);
   U1797 : NOR2_X1 port map( A1 => n8066, A2 => n7867, ZN => n4379);
   U1798 : BUF_X2 port map( A => n7047, Z => n7556);
   U1799 : BUF_X1 port map( A => n4561, Z => n5398);
   U1800 : BUF_X1 port map( A => n6705, Z => n4401);
   U1807 : INV_X1 port map( A => n7616, ZN => n4362);
   U1808 : NOR2_X1 port map( A1 => n8082, A2 => n4529, ZN => n8083);
   U1817 : OR2_X1 port map( A1 => n7368, A2 => n4450, ZN => n8123);
   U1818 : OR2_X1 port map( A1 => n7370, A2 => n7371, ZN => n7597);
   U1819 : BUF_X1 port map( A => n6668, Z => n4476);
   U1820 : CLKBUF_X1 port map( A => n4413, Z => n6557);
   U1821 : XNOR2_X1 port map( A => n7353, B => n7385, ZN => n8181);
   U1823 : XNOR2_X1 port map( A => n4378, B => n5830, ZN => n5571);
   U1828 : AOI22_X1 port map( A1 => n4396, A2 => n4395, B1 => n4925, B2 => 
                           n4924, ZN => n4929);
   U1833 : NAND2_X1 port map( A1 => n7971, A2 => n7800, ZN => n7801);
   U1834 : OR2_X1 port map( A1 => n6665, A2 => n6664, ZN => n4373);
   U1835 : AND2_X1 port map( A1 => n4909, A2 => n4910, ZN => n4398);
   U1836 : AND2_X1 port map( A1 => n5541, A2 => n5542, ZN => n5559);
   U1838 : INV_X1 port map( A => n8600, ZN => n6682);
   U1839 : XNOR2_X1 port map( A => n6027, B => n6206, ZN => n6522);
   U1840 : CLKBUF_X1 port map( A => n5179, Z => n4424);
   U1841 : CLKBUF_X1 port map( A => n5017, Z => n5018);
   U1842 : AND2_X1 port map( A1 => n4677, A2 => n4746, ZN => n4935);
   U1843 : NAND2_X1 port map( A1 => n4371, A2 => n4370, ZN => n5374);
   U1844 : OR2_X1 port map( A1 => n5453, A2 => n5452, ZN => n5580);
   U1845 : NOR2_X1 port map( A1 => n5977, A2 => n4385, ZN => n4384);
   U1846 : OR3_X1 port map( A1 => n8315, A2 => n8377, A3 => n8289, ZN => n8291)
                           ;
   U1847 : OR3_X1 port map( A1 => n8315, A2 => n2582, A3 => n8289, ZN => n8290)
                           ;
   U1848 : INV_X1 port map( A => n5972, ZN => n4385);
   U1850 : NAND2_X1 port map( A1 => n5183, A2 => n5182, ZN => n4370);
   U1852 : INV_X1 port map( A => n4403, ZN => n6419);
   U1854 : INV_X1 port map( A => n4836, ZN => n4865);
   U1858 : NAND4_X1 port map( A1 => n4837, A2 => n4841, A3 => n4844, A4 => 
                           n4898, ZN => n4836);
   U1860 : NAND2_X1 port map( A1 => n4821, A2 => n4820, ZN => n4898);
   U1861 : NAND2_X1 port map( A1 => n4390, A2 => n4391, ZN => n4389);
   U1864 : OAI21_X1 port map( B1 => n5994, B2 => n6165, A => n6164, ZN => n6162
                           );
   U1867 : INV_X1 port map( A => n6406, ZN => n4390);
   U1868 : XNOR2_X1 port map( A => n4814, B => n4841, ZN => n4837);
   U1871 : INV_X1 port map( A => n6405, ZN => n4391);
   U1872 : AND2_X1 port map( A1 => n4379, A2 => n7860, ZN => n8109);
   U1873 : AND2_X1 port map( A1 => n5897, A2 => n5896, ZN => n5952);
   U1874 : INV_X1 port map( A => n5627, ZN => n5625);
   U1875 : MUX2_X1 port map( A => n4462, B => n7198, S => n8396, Z => n5478);
   U1877 : AND2_X1 port map( A1 => n8093, A2 => n7859, ZN => n7860);
   U1878 : OR2_X1 port map( A1 => n5618, A2 => n5619, ZN => n5627);
   U1879 : NAND2_X1 port map( A1 => n7095, A2 => n390, ZN => n4368);
   U1881 : CLKBUF_X1 port map( A => n5937, Z => n5748);
   U1883 : BUF_X1 port map( A => n6889, Z => n4489);
   U1885 : BUF_X1 port map( A => n4573, Z => n4975);
   U1888 : NAND2_X1 port map( A1 => n5142, A2 => n6705, ZN => n7415);
   U1892 : BUF_X1 port map( A => n4560, Z => n5397);
   U1896 : NAND2_X1 port map( A1 => n4727, A2 => n8002, ZN => n6388);
   U1897 : BUF_X1 port map( A => n4727, Z => n6264);
   U1898 : CLKBUF_X3 port map( A => n5508, Z => n6595);
   U1899 : NAND2_X1 port map( A1 => n5386, A2 => n6113, ZN => n6696);
   U1901 : CLKBUF_X1 port map( A => n6113, Z => n6234);
   U1904 : AND2_X1 port map( A1 => n8356, A2 => n366, ZN => n4364);
   U1906 : NOR2_X1 port map( A1 => n4363, A2 => n4362, ZN => n7628);
   U1907 : OAI21_X1 port map( B1 => n8152, B2 => n7617, A => n7615, ZN => n4363
                           );
   U1909 : INV_X1 port map( A => n6056, ZN => n4365);
   U1910 : OAI21_X1 port map( B1 => n4366, B2 => n4367, A => n8128, ZN => n8139
                           );
   U1911 : OAI21_X1 port map( B1 => n8125, B2 => n4399, A => n8123, ZN => n4366
                           );
   U1912 : INV_X1 port map( A => n8124, ZN => n4367);
   U1914 : NAND2_X1 port map( A1 => n4368, A2 => n4369, ZN => n5868);
   U1915 : NAND2_X1 port map( A1 => n7096, A2 => n8352, ZN => n4369);
   U1916 : OAI21_X1 port map( B1 => n5183, B2 => n5182, A => n5181, ZN => n4371
                           );
   U1917 : NAND2_X1 port map( A1 => n5179, A2 => n5178, ZN => n5177);
   U1918 : XNOR2_X1 port map( A => n4372, B => n5183, ZN => n5179);
   U1919 : XNOR2_X1 port map( A => n5181, B => n5182, ZN => n4372);
   U1920 : AND3_X1 port map( A1 => n4373, A2 => n6663, A3 => n6662, ZN => n6680
                           );
   U1921 : NAND3_X1 port map( A1 => n8224, A2 => n8225, A3 => n4374, ZN => 
                           I2_dtemp_43_port);
   U1922 : NOR2_X1 port map( A1 => n4359, A2 => n4357, ZN => n4374);
   U1923 : NAND2_X1 port map( A1 => n6425, A2 => n8429, ZN => n4375);
   U1924 : OR2_X1 port map( A1 => n5706, A2 => n5705, ZN => n4377);
   U1925 : NAND2_X1 port map( A1 => n4478, A2 => n4691, ZN => n4587);
   U1926 : NAND2_X1 port map( A1 => n4557, A2 => n4558, ZN => n4691);
   U1929 : INV_X1 port map( A => n6162, ZN => n6172);
   U1932 : NAND2_X1 port map( A1 => n4377, A2 => n5704, ZN => n6071);
   U1934 : NOR2_X2 port map( A1 => n8261, A2 => n8260, ZN => n8259);
   U1935 : NAND2_X1 port map( A1 => n4382, A2 => n4380, ZN => n6125);
   U1937 : NAND2_X1 port map( A1 => n4437, A2 => n373, ZN => n4382);
   U1938 : NAND3_X1 port map( A1 => n5975, A2 => n5976, A3 => n4383, ZN => 
                           n6076);
   U1939 : NAND2_X1 port map( A1 => n5974, A2 => n4384, ZN => n4383);
   U1940 : NAND3_X1 port map( A1 => n4389, A2 => n4387, A3 => n4386, ZN => 
                           n4403);
   U1941 : NAND3_X1 port map( A1 => n4392, A2 => n6378, A3 => n4391, ZN => 
                           n4386);
   U1942 : NAND3_X1 port map( A1 => n6407, A2 => n6406, A3 => n6405, ZN => 
                           n4387);
   U1943 : INV_X1 port map( A => n6380, ZN => n4392);
   U1944 : NAND2_X1 port map( A1 => n4393, A2 => n4986, ZN => n4988);
   U1945 : NAND2_X1 port map( A1 => n4987, A2 => n4393, ZN => n4738);
   U1946 : NAND2_X1 port map( A1 => n4734, A2 => n4733, ZN => n4393);
   U1950 : INV_X1 port map( A => n4837, ZN => n4900);
   U1951 : OR2_X1 port map( A1 => n4923, A2 => n4922, ZN => n4395);
   U1952 : NAND3_X1 port map( A1 => n4398, A2 => n4911, A3 => n4397, ZN => 
                           n4396);
   U1953 : NAND2_X1 port map( A1 => n4922, A2 => n4923, ZN => n4397);
   U1954 : OR2_X1 port map( A1 => n4568, A2 => n4569, ZN => n4649);
   U1957 : NOR2_X1 port map( A1 => n8098, A2 => n7492, ZN => n7727);
   U1958 : XNOR2_X1 port map( A => n4420, B => n5171, ZN => n5174);
   U1959 : AND2_X1 port map( A1 => n8037, A2 => n8036, ZN => n8031);
   U1962 : AND2_X1 port map( A1 => n5114, A2 => n5113, ZN => n4405);
   U1963 : XOR2_X1 port map( A => n6600, B => n6599, Z => n4406);
   U1964 : NAND2_X1 port map( A1 => n5155, A2 => n5154, ZN => n4407);
   U1965 : OR2_X1 port map( A1 => n6877, A2 => n6878, ZN => n4408);
   U1966 : XOR2_X1 port map( A => n4407, B => n5156, Z => n4409);
   U1970 : INV_X1 port map( A => n8340, ZN => n4411);
   U1972 : XNOR2_X1 port map( A => n6533, B => n6532, ZN => n4413);
   U1973 : NAND2_X1 port map( A1 => n8204, A2 => n8209, ZN => n4414);
   U1974 : AND2_X1 port map( A1 => n5607, A2 => n5606, ZN => n4415);
   U1976 : NAND2_X1 port map( A1 => n4459, A2 => n7495, ZN => n4418);
   U1978 : NOR2_X1 port map( A1 => n6223, A2 => n6224, ZN => n7855);
   U1979 : XNOR2_X1 port map( A => n5173, B => n5172, ZN => n4420);
   U1980 : XNOR2_X1 port map( A => n4422, B => n6931, ZN => n4421);
   U1981 : XOR2_X1 port map( A => n6734, B => n4416, Z => n4422);
   U1983 : INV_X1 port map( A => n4430, ZN => n5407);
   U1984 : NAND2_X1 port map( A1 => n6640, A2 => n6641, ZN => n4425);
   U1985 : OR2_X1 port map( A1 => n8526, A2 => n7618, ZN => n4428);
   U1987 : XNOR2_X1 port map( A => n393, B => n370, ZN => n4430);
   U1988 : AND2_X1 port map( A1 => n6527, A2 => n6526, ZN => n4431);
   U1989 : NOR2_X1 port map( A1 => n6878, A2 => n6877, ZN => n6895);
   U1990 : NAND3_X1 port map( A1 => n7593, A2 => n7592, A3 => n4358, ZN => 
                           I2_dtemp_42_port);
   U1991 : OR2_X1 port map( A1 => n7485, A2 => n7486, ZN => n4432);
   U1992 : OR2_X1 port map( A1 => n7486, A2 => n7485, ZN => n7737);
   U1993 : NAND2_X1 port map( A1 => n6093, A2 => n6091, ZN => n4433);
   U1994 : XOR2_X1 port map( A => n6037, B => n6036, Z => n4434);
   U1995 : OR2_X1 port map( A1 => n6310, A2 => n6311, ZN => n6330);
   U1996 : AND2_X1 port map( A1 => n6802, A2 => n6801, ZN => n4435);
   U1997 : AND2_X1 port map( A1 => n6636, A2 => n6635, ZN => n4436);
   U2000 : AND3_X1 port map( A1 => n8527, A2 => n7624, A3 => n4532, ZN => n4438
                           );
   U2001 : NAND2_X1 port map( A1 => n6694, A2 => n4439, ZN => n6844);
   U2002 : AND2_X1 port map( A1 => n6693, A2 => n6843, ZN => n4439);
   U2003 : NAND2_X1 port map( A1 => n8468, A2 => n6844, ZN => n4440);
   U2006 : AND2_X1 port map( A1 => n7378, A2 => n7607, ZN => n4441);
   U2007 : OR2_X1 port map( A1 => n7174, A2 => n7173, ZN => n4442);
   U2013 : OAI21_X1 port map( B1 => n8597, B2 => n6087, A => n6086, ZN => n4447
                           );
   U2014 : OAI21_X1 port map( B1 => n8517, B2 => n6087, A => n6086, ZN => n8204
                           );
   U2015 : OAI211_X1 port map( C1 => n6991, C2 => n6990, A => n6989, B => n8464
                           , ZN => n4448);
   U2016 : BUF_X1 port map( A => n7983, Z => n4449);
   U2017 : BUF_X2 port map( A => n389, Z => n8002);
   U2018 : NAND2_X1 port map( A1 => n7095, A2 => n356, ZN => n4509);
   U2020 : INV_X1 port map( A => n387, ZN => n6113);
   U2022 : INV_X1 port map( A => n5008, ZN => n5009);
   U2023 : NAND2_X1 port map( A1 => n6113, A2 => n8364, ZN => n5937);
   U2024 : OR2_X1 port map( A1 => n6895, A2 => n6896, ZN => n7060);
   U2026 : NAND2_X1 port map( A1 => n6358, A2 => n6357, ZN => n6587);
   U2027 : NAND2_X1 port map( A1 => n6588, A2 => n6590, ZN => n6592);
   U2028 : NAND2_X1 port map( A1 => n7060, A2 => n4519, ZN => n7154);
   U2029 : NAND2_X1 port map( A1 => n7061, A2 => n7062, ZN => n4519);
   U2030 : NAND2_X1 port map( A1 => n5564, A2 => n5563, ZN => n5573);
   U2031 : XNOR2_X1 port map( A => n5559, B => n5558, ZN => n5562);
   U2032 : OR2_X1 port map( A1 => n4979, A2 => n4978, ZN => n5112);
   U2033 : NOR2_X1 port map( A1 => n7298, A2 => n7297, ZN => n7302);
   U2035 : INV_X1 port map( A => n7032, ZN => n7035);
   U2038 : OAI21_X1 port map( B1 => n6715, B2 => n379, A => n4454, ZN => n4453)
                           ;
   U2039 : NAND2_X1 port map( A1 => n5872, A2 => n379, ZN => n4454);
   U2040 : NAND2_X1 port map( A1 => n7119, A2 => n7118, ZN => n7152);
   U2041 : INV_X1 port map( A => n7062, ZN => n6898);
   U2042 : AND2_X1 port map( A1 => n6609, A2 => n8504, ZN => n6610);
   U2043 : INV_X1 port map( A => n6613, ZN => n6615);
   U2045 : AND2_X1 port map( A1 => n5863, A2 => n5862, ZN => n6175);
   U2047 : OAI22_X1 port map( A1 => n4518, A2 => n6587, B1 => n6592, B2 => 
                           n6589, ZN => n6734);
   U2048 : AOI21_X1 port map( B1 => n6588, B2 => n6590, A => n6591, ZN => n4518
                           );
   U2051 : XNOR2_X1 port map( A => n5264, B => n5178, ZN => n5153);
   U2053 : AND3_X1 port map( A1 => n7640, A2 => n7481, A3 => n7482, ZN => n7723
                           );
   U2054 : INV_X1 port map( A => n8131, ZN => n7594);
   U2055 : INV_X1 port map( A => n7154, ZN => n7153);
   U2056 : OR2_X1 port map( A1 => n6602, A2 => n6948, ZN => n6601);
   U2058 : NOR2_X1 port map( A1 => n7801, A2 => n4525, ZN => n4524);
   U2059 : INV_X1 port map( A => n7805, ZN => n4525);
   U2060 : INV_X1 port map( A => n8080, ZN => n8082);
   U2061 : NAND2_X1 port map( A1 => n6804, A2 => n6803, ZN => n6997);
   U2062 : NAND2_X1 port map( A1 => n8478, A2 => n205, ZN => n6821);
   U2063 : AND2_X1 port map( A1 => n8370, A2 => n8395, ZN => n4538);
   U2064 : AND2_X1 port map( A1 => n5104, A2 => n5103, ZN => n5108);
   U2065 : OR2_X1 port map( A1 => n5353, A2 => n5351, ZN => n5350);
   U2067 : BUF_X1 port map( A => n392, Z => n5848);
   U2068 : INV_X1 port map( A => n6997, ZN => n7001);
   U2069 : NAND2_X1 port map( A1 => n8401, A2 => n8350, ZN => n6607);
   U2070 : NAND2_X1 port map( A1 => n6459, A2 => n6458, ZN => n6469);
   U2071 : MUX2_X1 port map( A => n7692, B => n7254, S => n8352, Z => n6459);
   U2073 : AND2_X1 port map( A1 => n5747, A2 => n8398, ZN => n5936);
   U2074 : OR2_X1 port map( A1 => n7100, A2 => n7099, ZN => n7180);
   U2075 : OR2_X1 port map( A1 => n7007, A2 => n7006, ZN => n7004);
   U2076 : INV_X1 port map( A => n6881, ZN => n4512);
   U2079 : INV_X1 port map( A => n6852, ZN => n6856);
   U2080 : OR2_X1 port map( A1 => n6757, A2 => n6753, ZN => n6758);
   U2082 : NAND2_X1 port map( A1 => n6040, A2 => n6039, ZN => n6044);
   U2083 : OR2_X1 port map( A1 => n6042, A2 => n6041, ZN => n6039);
   U2084 : OAI211_X1 port map( C1 => n7227, C2 => n386, A => n5647, B => n4530,
                           ZN => n5721);
   U2085 : NOR2_X1 port map( A1 => n5345, A2 => n5344, ZN => n5676);
   U2086 : NAND2_X1 port map( A1 => n5447, A2 => n4452, ZN => n5512);
   U2087 : INV_X1 port map( A => n4453, ZN => n4452);
   U2088 : NOR2_X1 port map( A1 => n5546, A2 => n5545, ZN => n5548);
   U2089 : OR2_X1 port map( A1 => n7262, A2 => n7261, ZN => n7350);
   U2090 : INV_X1 port map( A => n6174, ZN => n6177);
   U2091 : INV_X1 port map( A => n5771, ZN => n5522);
   U2092 : OR2_X1 port map( A1 => n5808, A2 => n5807, ZN => n6054);
   U2093 : CLKBUF_X1 port map( A => n7922, Z => n7924);
   U2094 : NAND2_X1 port map( A1 => n7188, A2 => n7187, ZN => n7355);
   U2095 : INV_X1 port map( A => n6970, ZN => n6925);
   U2096 : CLKBUF_X1 port map( A => n6962, Z => n6963);
   U2097 : XNOR2_X1 port map( A => n4511, B => n6647, ZN => n6660);
   U2098 : XNOR2_X1 port map( A => n6646, B => n6645, ZN => n4511);
   U2099 : INV_X1 port map( A => n6292, ZN => n4513);
   U2101 : INV_X1 port map( A => n6959, ZN => n6624);
   U2102 : NAND2_X1 port map( A1 => n6219, A2 => n6218, ZN => n6220);
   U2103 : NOR2_X1 port map( A1 => n6219, A2 => n6218, ZN => n6222);
   U2105 : NOR2_X1 port map( A1 => n4522, A2 => n4523, ZN => n8367);
   U2108 : AND2_X1 port map( A1 => n6780, A2 => n6779, ZN => n4450);
   U2109 : AOI22_X1 port map( A1 => n4456, A2 => n6936, B1 => n6935, B2 => 
                           n6934, ZN => n6971);
   U2110 : OR2_X1 port map( A1 => n8605, A2 => n7966, ZN => n4451);
   U2111 : AND2_X2 port map( A1 => n6817, A2 => n8368, ZN => n5872);
   U2112 : XOR2_X1 port map( A => n6772, B => n6771, Z => n4456);
   U2113 : XNOR2_X1 port map( A => n5246, B => n5333, ZN => n4457);
   U2115 : NAND2_X1 port map( A1 => n6608, A2 => n6607, ZN => n6611);
   U2116 : AND2_X1 port map( A1 => n5611, A2 => n5610, ZN => n4458);
   U2118 : XOR2_X1 port map( A => n391, B => n164, Z => n4727);
   U2119 : OR2_X1 port map( A1 => n5431, A2 => n5430, ZN => n4460);
   U2122 : AND2_X1 port map( A1 => n4484, A2 => n7165, ZN => n7162);
   U2123 : OAI21_X1 port map( B1 => n7771, B2 => n4381, A => n7033, ZN => n7034
                           );
   U2125 : XOR2_X1 port map( A => n5821, B => n8540, Z => n4464);
   U2126 : NAND2_X1 port map( A1 => n7009, A2 => n7008, ZN => n4465);
   U2128 : OR2_X1 port map( A1 => n8181, A2 => n8180, ZN => n7599);
   U2129 : XNOR2_X1 port map( A => n7267, B => n7349, ZN => n4467);
   U2130 : AND3_X1 port map( A1 => n8497, A2 => n5029, A3 => n5027, ZN => n4468
                           );
   U2131 : NAND2_X1 port map( A1 => n5516, A2 => n5550, ZN => n4469);
   U2132 : NAND2_X1 port map( A1 => n5516, A2 => n8570, ZN => n4470);
   U2133 : NAND2_X1 port map( A1 => n5550, A2 => n8570, ZN => n4471);
   U2135 : NAND2_X1 port map( A1 => n5104, A2 => n5103, ZN => n4472);
   U2136 : NAND2_X1 port map( A1 => n6694, A2 => n6693, ZN => n4473);
   U2137 : MUX2_X1 port map( A => n7120, B => n7121, S => n8328, Z => n4965);
   U2139 : NOR2_X1 port map( A1 => n6979, A2 => n6980, ZN => n4474);
   U2140 : NAND2_X1 port map( A1 => n6982, A2 => n6981, ZN => n4475);
   U2141 : NAND2_X1 port map( A1 => n7148, A2 => n7147, ZN => n7185);
   U2145 : OR2_X1 port map( A1 => n4558, A2 => n4557, ZN => n4478);
   U2146 : NAND2_X1 port map( A1 => n5020, A2 => n5019, ZN => n4479);
   U2147 : NAND2_X1 port map( A1 => n5020, A2 => n5018, ZN => n4480);
   U2148 : NAND2_X1 port map( A1 => n5019, A2 => n5018, ZN => n4481);
   U2149 : NAND3_X1 port map( A1 => n4479, A2 => n4480, A3 => n4481, ZN => 
                           n5175);
   U2150 : INV_X1 port map( A => n5016, ZN => n5019);
   U2151 : XNOR2_X1 port map( A => n5826, B => n5825, ZN => n8037);
   U2153 : AND2_X1 port map( A1 => n8484, A2 => n8073, ZN => n4482);
   U2154 : XNOR2_X1 port map( A => n367, B => n392, ZN => n4817);
   U2157 : AND2_X1 port map( A1 => n7068, A2 => n7067, ZN => n4484);
   U2158 : NAND2_X1 port map( A1 => n7367, A2 => n7366, ZN => n4485);
   U2159 : NAND2_X1 port map( A1 => n6785, A2 => n6784, ZN => n4486);
   U2162 : XNOR2_X1 port map( A => n8506, B => A_SIG_10_port, ZN => n4491);
   U2163 : NAND2_X1 port map( A1 => n4658, A2 => n5883, ZN => n6889);
   U2164 : XOR2_X1 port map( A => n6543, B => n6558, Z => n4492);
   U2165 : XNOR2_X1 port map( A => n6288, B => n4513, ZN => n6536);
   U2166 : NAND2_X1 port map( A1 => n6062, A2 => n6063, ZN => n4493);
   U2167 : NAND2_X1 port map( A1 => n6062, A2 => n8467, ZN => n4494);
   U2168 : NAND2_X1 port map( A1 => n6063, A2 => n8467, ZN => n4495);
   U2169 : NAND3_X1 port map( A1 => n4493, A2 => n4494, A3 => n4495, ZN => 
                           n8050);
   U2170 : XOR2_X1 port map( A => n5963, B => n8557, Z => n4496);
   U2171 : XOR2_X1 port map( A => n5953, B => n5952, Z => n4497);
   U2172 : OR2_X1 port map( A1 => n4448, A2 => n7477, ZN => n4498);
   U2173 : XNOR2_X1 port map( A => n7237, B => n7085, ZN => n7104);
   U2174 : INV_X2 port map( A => n5794, ZN => n6102);
   U2176 : XNOR2_X1 port map( A => n8569, B => n6052, ZN => n6221);
   U2177 : AOI21_X1 port map( B1 => n4957, B2 => n4956, A => n4955, ZN => n4499
                           );
   U2178 : AND2_X1 port map( A1 => n4498, A2 => n8157, ZN => n4500);
   U2179 : OR2_X1 port map( A1 => n4734, A2 => n4733, ZN => n4987);
   U2180 : OR2_X1 port map( A1 => n8077, A2 => n4444, ZN => n7623);
   U2181 : OR2_X1 port map( A1 => n7642, A2 => n7633, ZN => n4501);
   U2182 : OR2_X1 port map( A1 => n4501, A2 => n7956, ZN => n7649);
   U2184 : AOI21_X1 port map( B1 => n6906, B2 => n6905, A => n6904, ZN => n7064
                           );
   U2185 : AOI21_X1 port map( B1 => n6905, B2 => n6903, A => n6906, ZN => n4515
                           );
   U2186 : OAI211_X1 port map( C1 => n4399, C2 => n8125, A => n8124, B => n8123
                           , ZN => n4503);
   U2187 : XOR2_X1 port map( A => n5554, B => n5555, Z => n4504);
   U2188 : AND2_X1 port map( A1 => n7972, A2 => n4524, ZN => n4523);
   U2189 : NAND2_X1 port map( A1 => n5623, A2 => n5622, ZN => n5626);
   U2190 : NOR2_X1 port map( A1 => n5251, A2 => n5252, ZN => n4506);
   U2191 : NAND2_X1 port map( A1 => n5166, A2 => n5165, ZN => n5253);
   U2192 : XNOR2_X1 port map( A => n4507, B => n5583, ZN => n5452);
   U2193 : XNOR2_X1 port map( A => n5584, B => n5586, ZN => n4507);
   U2194 : NOR2_X1 port map( A1 => n7723, A2 => n7728, ZN => n7724);
   U2195 : NAND3_X1 port map( A1 => n7964, A2 => n7965, A3 => n4451, ZN => 
                           I2_dtemp_40_port);
   U2196 : NAND2_X1 port map( A1 => n8131, A2 => n8103, ZN => n7602);
   U2198 : NOR2_X1 port map( A1 => n6807, A2 => n4508, ZN => n6810);
   U2199 : NAND2_X1 port map( A1 => n4510, A2 => n4509, ZN => n4508);
   U2200 : NAND2_X1 port map( A1 => n7096, A2 => n8326, ZN => n4510);
   U2201 : MUX2_X1 port map( A => n7121, B => n7120, S => n8423, Z => n6815);
   U2202 : MUX2_X1 port map( A => n7121, B => n7120, S => n6606, Z => n5068);
   U2203 : MUX2_X1 port map( A => n7121, B => n7120, S => n359, Z => n6307);
   U2204 : MUX2_X1 port map( A => n7121, B => n7120, S => n204, Z => n5650);
   U2205 : MUX2_X1 port map( A => n7121, B => n7120, S => n379, Z => n5945);
   U2206 : INV_X1 port map( A => n4515, ZN => n4516);
   U2207 : NAND3_X1 port map( A1 => n4517, A2 => n6871, A3 => n4516, ZN => 
                           n6942);
   U2208 : NAND3_X1 port map( A1 => n6905, A2 => n6906, A3 => n6903, ZN => 
                           n4517);
   U2209 : NAND2_X1 port map( A1 => n6941, A2 => n6942, ZN => n6944);
   U2210 : NOR2_X1 port map( A1 => n8526, A2 => n7618, ZN => n8146);
   U2211 : NOR2_X1 port map( A1 => n8123, A2 => n7594, ZN => n7618);
   U2213 : NAND2_X1 port map( A1 => n7983, A2 => n7989, ZN => n7972);
   U2214 : OAI21_X1 port map( B1 => n5562, B2 => n5561, A => n5560, ZN => n5564
                           );
   U2216 : OR2_X1 port map( A1 => n7626, A2 => n8144, ZN => n7627);
   U2217 : BUF_X1 port map( A => n8152, Z => n8184);
   U2219 : NAND2_X1 port map( A1 => n4693, A2 => n4478, ZN => n5016);
   U2221 : NAND2_X1 port map( A1 => n6290, A2 => n6289, ZN => n6544);
   U2222 : OR2_X1 port map( A1 => n7059, A2 => n7058, ZN => n7156);
   U2224 : XNOR2_X1 port map( A => n7239, B => n7235, ZN => n7085);
   U2227 : XNOR2_X1 port map( A => A_SIG_16_port, B => n384, ZN => n5142);
   U2228 : OR2_X1 port map( A1 => n7478, A2 => n7477, ZN => n8149);
   U2229 : NAND2_X1 port map( A1 => n5407, A2 => n8503, ZN => n7086);
   U2230 : OAI21_X1 port map( B1 => n6538, B2 => n6534, A => n6536, ZN => n6290
                           );
   U2231 : XNOR2_X1 port map( A => n6266, B => n6443, ZN => n6538);
   U2232 : NAND2_X1 port map( A1 => n5508, A2 => n6343, ZN => n5866);
   U2233 : OAI22_X1 port map( A1 => n8004, A2 => n8329, B1 => n8003, B2 => n363
                           , ZN => n5865);
   U2234 : OR2_X1 port map( A1 => n7323, A2 => n395, ZN => n4526);
   U2236 : OR2_X1 port map( A1 => n8279, A2 => SIG_in_26_port, ZN => n4527);
   U2237 : AND2_X1 port map( A1 => n6264, A2 => n5864, ZN => n4528);
   U2238 : AND3_X1 port map( A1 => n6564, A2 => n6563, A3 => n8081, ZN => n4529
                           );
   U2239 : OR2_X1 port map( A1 => n7439, A2 => n8328, ZN => n4530);
   U2240 : AND2_X1 port map( A1 => n7808, A2 => n7807, ZN => n4531);
   U2241 : AND4_X1 port map( A1 => n7623, A2 => n8541, A3 => n7734, A4 => n7621
                           , ZN => n4532);
   U2243 : BUF_X1 port map( A => n5030, Z => n7121);
   U2244 : AND3_X1 port map( A1 => n8586, A2 => n8075, A3 => n8490, ZN => n4533
                           );
   U2245 : CLKBUF_X1 port map( A => n5898, Z => n4867);
   U2246 : AOI21_X1 port map( B1 => n4849, B2 => n4903, A => n4904, ZN => n4866
                           );
   U2247 : INV_X1 port map( A => n5120, ZN => n4960);
   U2248 : OR2_X1 port map( A1 => n6688, A2 => n360, ZN => n6690);
   U2249 : AOI21_X1 port map( B1 => n4957, B2 => n4956, A => n4955, ZN => n5116
                           );
   U2252 : BUF_X1 port map( A => n383, Z => n5273);
   U2253 : NAND2_X1 port map( A1 => n4697, A2 => n4696, ZN => n5008);
   U2254 : NAND2_X1 port map( A1 => n7087, A2 => n377, ZN => n7088);
   U2256 : INV_X1 port map( A => n6839, ZN => n6840);
   U2257 : OAI22_X1 port map( A1 => n7392, A2 => B_SIG_8_port, B1 => n8362, B2 
                           => n7253, ZN => n6614);
   U2258 : NAND2_X1 port map( A1 => n4997, A2 => n384, ZN => n6688);
   U2259 : OR2_X1 port map( A1 => n5351, A2 => n5352, ZN => n5347);
   U2260 : OAI211_X1 port map( C1 => n7324, C2 => n8393, A => n5043, B => n4526
                           , ZN => n5047);
   U2261 : NAND2_X1 port map( A1 => n5148, A2 => n4356, ZN => n5150);
   U2262 : OR2_X1 port map( A1 => n4984, A2 => n4985, ZN => n5160);
   U2264 : OR2_X1 port map( A1 => n7015, A2 => n7128, ZN => n7146);
   U2265 : INV_X1 port map( A => n8458, ZN => n6854);
   U2266 : NAND2_X1 port map( A1 => n6717, A2 => n6716, ZN => n6852);
   U2267 : NOR2_X1 port map( A1 => n6615, A2 => n6614, ZN => n6616);
   U2268 : OR2_X1 port map( A1 => n5677, A2 => n5674, ZN => n5491);
   U2269 : NAND2_X1 port map( A1 => n5150, A2 => n8537, ZN => n5206);
   U2270 : OR2_X1 port map( A1 => n4926, A2 => intadd_33_n1, ZN => n4772);
   U2271 : INV_X1 port map( A => n8399, ZN => n5777);
   U2272 : OR2_X1 port map( A1 => n7239, A2 => n7238, ZN => n7236);
   U2273 : NAND2_X1 port map( A1 => n6783, A2 => n6782, ZN => n7021);
   U2274 : XNOR2_X1 port map( A => n6281, B => n6280, ZN => n6108);
   U2275 : INV_X1 port map( A => n5206, ZN => n5151);
   U2276 : NAND2_X1 port map( A1 => n6042, A2 => n6041, ZN => n6043);
   U2277 : NOR2_X1 port map( A1 => n7174, A2 => n7173, ZN => n7177);
   U2278 : INV_X1 port map( A => n7185, ZN => n7149);
   U2279 : OR2_X1 port map( A1 => n4440, A2 => n6867, ZN => n6905);
   U2280 : NOR2_X1 port map( A1 => n8587, A2 => n8599, ZN => n6932);
   U2281 : INV_X1 port map( A => n6496, ZN => n6332);
   U2282 : XNOR2_X1 port map( A => n6108, B => n6279, ZN => n6268);
   U2283 : NOR2_X1 port map( A1 => n7269, A2 => n7242, ZN => n7248);
   U2284 : OR2_X1 port map( A1 => n7457, A2 => n7458, ZN => n7460);
   U2285 : AND2_X1 port map( A1 => n7599, A2 => n8175, ZN => n7381);
   U2286 : OR2_X1 port map( A1 => n5507, A2 => n5506, ZN => n5526);
   U2287 : NAND2_X1 port map( A1 => n6044, A2 => n6043, ZN => n6050);
   U2288 : AND2_X1 port map( A1 => n4443, A2 => n7189, ZN => n7194);
   U2289 : XNOR2_X1 port map( A => n6722, B => n6623, ZN => n6958);
   U2290 : XNOR2_X1 port map( A => n5871, B => n6137, ZN => n5910);
   U2291 : NAND2_X1 port map( A1 => n6538, A2 => n6534, ZN => n6289);
   U2292 : NAND2_X1 port map( A1 => n5639, A2 => n5636, ZN => n5771);
   U2293 : INV_X1 port map( A => n5557, ZN => n5558);
   U2294 : AND2_X1 port map( A1 => n7988, A2 => n7734, ZN => n7736);
   U2295 : NAND2_X1 port map( A1 => n6049, A2 => n6050, ZN => n6057);
   U2296 : XNOR2_X1 port map( A => n4424, B => n5153, ZN => n5265);
   U2297 : NAND2_X1 port map( A1 => n7286, A2 => n7285, ZN => n7287);
   U2298 : NAND2_X1 port map( A1 => n5562, A2 => n5561, ZN => n5563);
   U2299 : NAND2_X1 port map( A1 => n7288, A2 => n7287, ZN => n7373);
   U2302 : OAI21_X1 port map( B1 => n6778, B2 => n6777, A => n8545, ZN => n6780
                           );
   U2303 : OAI21_X1 port map( B1 => n6222, B2 => n6221, A => n6220, ZN => n6224
                           );
   U2304 : AND2_X1 port map( A1 => n8127, A2 => n8130, ZN => n8128);
   n8317 <= '1';
   n8318 <= '0';
   U2312 : NOR2_X1 port map( A1 => n4817, A2 => n5879, ZN => n4573);
   U2313 : INV_X1 port map( A => n4573, ZN => n5844);
   U2314 : NOR2_X1 port map( A1 => n4817, A2 => n8397, ZN => n4574);
   U2315 : INV_X1 port map( A => n4574, ZN => n5845);
   U2316 : MUX2_X1 port map( A => n5844, B => n5845, S => B_SIG_9_port, Z => 
                           n4535);
   U2317 : NAND2_X1 port map( A1 => n367, A2 => n392, ZN => n4810);
   U2318 : BUF_X2 port map( A => n391, Z => n4809);
   U2320 : INV_X1 port map( A => n8553, ZN => n5878);
   U2321 : NOR2_X1 port map( A1 => n367, A2 => n392, ZN => n4808);
   U2322 : BUF_X2 port map( A => B_SIG_8_port, Z => n6109);
   U2323 : MUX2_X1 port map( A => n6103, B => n6102, S => n6109, Z => n4534);
   U2324 : NAND2_X1 port map( A1 => n4535, A2 => n4534, ZN => n4718);
   U2325 : XNOR2_X1 port map( A => n366, B => n385, ZN => n4885);
   U2327 : INV_X1 port map( A => n5396, ZN => n5898);
   U2328 : NAND2_X1 port map( A1 => n5898, A2 => n8392, ZN => n4537);
   U2329 : NOR2_X1 port map( A1 => n4885, A2 => n5848, ZN => n4559);
   U2331 : NAND2_X1 port map( A1 => n6249, A2 => n379, ZN => n4536);
   U2332 : NAND2_X1 port map( A1 => n4537, A2 => n4536, ZN => n4540);
   U2333 : BUF_X2 port map( A => n385, Z => n6259);
   U2335 : MUX2_X1 port map( A => n6126, B => n6248, S => n204, Z => n4539);
   U2336 : NAND2_X1 port map( A1 => n4540, A2 => n4539, ZN => n4719);
   U2337 : XNOR2_X1 port map( A => n4719, B => n4718, ZN => n4543);
   U2338 : XNOR2_X1 port map( A => A_SIG_8_port, B => n389, ZN => n5051);
   U2339 : NAND2_X1 port map( A1 => n5051, A2 => n6244, ZN => n6714);
   U2342 : MUX2_X1 port map( A => n6714, B => n6888, S => n6606, Z => n4542);
   U2343 : NAND3_X1 port map( A1 => A_SIG_8_port, A2 => n388, A3 => n8355, ZN 
                           => n6819);
   U2344 : BUF_X2 port map( A => n6819, Z => n6715);
   U2345 : NOR2_X1 port map( A1 => n8355, A2 => n388, ZN => n6817);
   U2346 : MUX2_X1 port map( A => n6715, B => n6887, S => n8324, Z => n4541);
   U2347 : AND2_X1 port map( A1 => n4542, A2 => n4541, ZN => n4723);
   U2348 : XNOR2_X1 port map( A => n4543, B => n4723, ZN => n4558);
   U2351 : NAND2_X1 port map( A1 => n4658, A2 => n8340, ZN => n4632);
   U2352 : MUX2_X1 port map( A => n4490, B => n8577, S => n386, Z => n4546);
   U2355 : NOR2_X1 port map( A1 => n8338, A2 => n382, ZN => n4544);
   U2357 : MUX2_X1 port map( A => n4607, B => n8595, S => n381, Z => n4545);
   U2358 : NAND2_X1 port map( A1 => n4546, A2 => n4545, ZN => n4737);
   U2359 : INV_X1 port map( A => n4737, ZN => n4556);
   U2361 : NAND3_X1 port map( A1 => n8403, A2 => n4411, A3 => n369, ZN => n4963
                           );
   U2363 : XNOR2_X1 port map( A => n8360, B => n382, ZN => n4962);
   U2364 : BUF_X1 port map( A => n8514, Z => n5307);
   U2365 : XNOR2_X1 port map( A => n4961, B => n8393, ZN => n4548);
   U2366 : NAND2_X1 port map( A1 => n5307, A2 => n4548, ZN => n4549);
   U2368 : MUX2_X1 port map( A => n7946, B => n7947, S => n356, Z => n4552);
   U2369 : NAND2_X1 port map( A1 => n8395, A2 => mult_x_19_n4, ZN => n7949);
   U2370 : INV_X2 port map( A => n7949, ZN => n5781);
   U2371 : NAND2_X1 port map( A1 => n5781, A2 => n373, ZN => n4551);
   U2372 : AND2_X1 port map( A1 => n4552, A2 => n4551, ZN => n4553);
   U2373 : NAND2_X1 port map( A1 => n8462, A2 => n4553, ZN => n4736);
   U2374 : NAND2_X1 port map( A1 => n4736, A2 => n4455, ZN => n4555);
   U2375 : XNOR2_X1 port map( A => n4555, B => n4556, ZN => n4557);
   U2376 : MUX2_X1 port map( A => n5395, B => n8488, S => B_SIG_9_port, Z => 
                           n4563);
   U2377 : MUX2_X1 port map( A => n5397, B => n5398, S => n7945, Z => n4562);
   U2378 : NOR2_X1 port map( A1 => n4563, A2 => n4562, ZN => n4568);
   U2379 : INV_X1 port map( A => n7051, ZN => n4565);
   U2380 : INV_X1 port map( A => n8595, ZN => n4564);
   U2381 : AOI21_X1 port map( B1 => n4565, B2 => n2638, A => n4564, ZN => n4569
                           );
   U2382 : NAND2_X1 port map( A1 => n4568, A2 => n4569, ZN => n4650);
   U2383 : MUX2_X1 port map( A => n6714, B => n6888, S => n386, Z => n4567);
   U2384 : MUX2_X1 port map( A => n6715, B => n6887, S => n381, Z => n4566);
   U2385 : NAND2_X1 port map( A1 => n4567, A2 => n4566, ZN => n4651);
   U2386 : NAND2_X1 port map( A1 => n4650, A2 => n4651, ZN => n4570);
   U2387 : NAND2_X1 port map( A1 => n4570, A2 => n4649, ZN => n4681);
   U2388 : NAND2_X2 port map( A1 => n4727, A2 => n8538, ZN => n6740);
   U2389 : MUX2_X1 port map( A => n8445, B => n6740, S => n376, Z => n4583);
   U2391 : MUX2_X1 port map( A => n7946, B => n7947, S => n379, Z => n4572);
   U2392 : NAND2_X1 port map( A1 => n5781, A2 => n204, ZN => n4571);
   U2393 : NAND2_X1 port map( A1 => n4572, A2 => n4571, ZN => n4579);
   U2394 : INV_X1 port map( A => n4579, ZN => n4630);
   U2395 : BUF_X1 port map( A => n4574, Z => n8012);
   U2396 : MUX2_X1 port map( A => n4975, B => n8012, S => n6109, Z => n4576);
   U2397 : MUX2_X1 port map( A => n8455, B => n8553, S => n362, Z => n4575);
   U2398 : NOR2_X1 port map( A1 => n4576, A2 => n4575, ZN => n4578);
   U2399 : INV_X1 port map( A => n8434, ZN => n5034);
   U2402 : INV_X1 port map( A => n8459, ZN => n5033);
   U2403 : MUX2_X1 port map( A => n5034, B => n5033, S => n8324, Z => n4581);
   U2404 : NAND2_X1 port map( A1 => n4581, A2 => n4579, ZN => n4577);
   U2405 : OAI211_X1 port map( C1 => n4583, C2 => n4630, A => n4578, B => n4577
                           , ZN => n4678);
   U2406 : NAND2_X1 port map( A1 => n4681, A2 => n4678, ZN => n4585);
   U2407 : INV_X1 port map( A => n4578, ZN => n4580);
   U2408 : AND2_X1 port map( A1 => n4580, A2 => n4579, ZN => n4584);
   U2409 : INV_X1 port map( A => n4581, ZN => n4582);
   U2410 : NAND2_X1 port map( A1 => n4583, A2 => n4582, ZN => n4631);
   U2411 : NAND2_X1 port map( A1 => n4584, A2 => n4631, ZN => n4679);
   U2412 : NAND2_X1 port map( A1 => n4585, A2 => n4679, ZN => n4690);
   U2413 : INV_X1 port map( A => n4690, ZN => n4586);
   U2414 : XNOR2_X1 port map( A => n4587, B => n4586, ZN => n4618);
   U2415 : NAND2_X1 port map( A1 => n4360, A2 => n7122, ZN => n7230);
   U2416 : NAND2_X1 port map( A1 => n7122, A2 => n8354, ZN => n4588);
   U2417 : AND2_X1 port map( A1 => n7230, A2 => n4588, ZN => n5006);
   U2418 : INV_X1 port map( A => n5006, ZN => n4592);
   U2419 : MUX2_X1 port map( A => n8445, B => n6740, S => n362, Z => n4695);
   U2420 : MUX2_X1 port map( A => n8459, B => n8434, S => n8352, Z => n4694);
   U2421 : NAND3_X1 port map( A1 => n4695, A2 => n4592, A3 => n4694, ZN => 
                           n4591);
   U2422 : INV_X1 port map( A => n4694, ZN => n4589);
   U2423 : NAND2_X1 port map( A1 => n5006, A2 => n4589, ZN => n4590);
   U2424 : OAI211_X1 port map( C1 => n4592, C2 => n4695, A => n4591, B => n4590
                           , ZN => n4603);
   U2425 : MUX2_X1 port map( A => n7946, B => n7947, S => n373, Z => n4594);
   U2426 : NAND2_X1 port map( A1 => n5781, A2 => n379, ZN => n4593);
   U2427 : NAND2_X1 port map( A1 => n4594, A2 => n4593, ZN => n4627);
   U2428 : INV_X1 port map( A => n5307, ZN => n4595);
   U2429 : NOR2_X1 port map( A1 => n4595, A2 => n2638, ZN => n4598);
   U2430 : NAND2_X1 port map( A1 => n4627, A2 => n4598, ZN => n4596);
   U2431 : MUX2_X1 port map( A => n8459, B => n8434, S => n8401, Z => n4624);
   U2432 : AND2_X1 port map( A1 => n4596, A2 => n4624, ZN => n4597);
   U2433 : MUX2_X1 port map( A => n8445, B => n6740, S => n8564, Z => n4625);
   U2434 : NAND2_X1 port map( A1 => n4597, A2 => n4625, ZN => n4601);
   U2435 : INV_X1 port map( A => n4627, ZN => n4599);
   U2436 : INV_X1 port map( A => n4598, ZN => n4626);
   U2437 : NAND2_X1 port map( A1 => n4599, A2 => n4626, ZN => n4600);
   U2438 : NAND2_X1 port map( A1 => n4601, A2 => n4600, ZN => n4602);
   U2439 : NOR2_X1 port map( A1 => n4603, A2 => n4602, ZN => n4741);
   U2440 : INV_X1 port map( A => n4741, ZN => n4604);
   U2441 : NAND2_X1 port map( A1 => n4603, A2 => n4602, ZN => n4739);
   U2442 : NAND2_X1 port map( A1 => n4604, A2 => n4739, ZN => n4616);
   U2443 : MUX2_X1 port map( A => n6714, B => n6888, S => n8324, Z => n4606);
   U2444 : INV_X1 port map( A => n5872, ZN => n6243);
   U2445 : MUX2_X1 port map( A => n6715, B => n6887, S => n386, Z => n4605);
   U2447 : MUX2_X1 port map( A => n4490, B => n7051, S => n381, Z => n4609);
   U2449 : MUX2_X1 port map( A => n4607, B => n8595, S => n395, Z => n4608);
   U2450 : NAND2_X1 port map( A1 => n4609, A2 => n4608, ZN => n4612);
   U2451 : MUX2_X1 port map( A => n5898, B => n6249, S => n204, Z => n4611);
   U2452 : MUX2_X1 port map( A => n8454, B => n8516, S => n8327, Z => n4610);
   U2453 : NAND2_X1 port map( A1 => n4611, A2 => n4610, ZN => n4620);
   U2454 : NAND2_X1 port map( A1 => n4612, A2 => n4620, ZN => n4614);
   U2455 : INV_X1 port map( A => n4612, ZN => n4622);
   U2456 : INV_X1 port map( A => n4620, ZN => n4613);
   U2457 : AOI22_X1 port map( A1 => n4619, A2 => n4614, B1 => n4622, B2 => 
                           n4613, ZN => n4740);
   U2458 : INV_X1 port map( A => n4740, ZN => n4615);
   U2459 : XNOR2_X1 port map( A => n4616, B => n4615, ZN => n4617);
   U2460 : NAND2_X1 port map( A1 => n4618, A2 => n4617, ZN => n4687);
   U2461 : NAND2_X1 port map( A1 => n4689, A2 => n4687, ZN => n4648);
   U2463 : XNOR2_X1 port map( A => n4621, B => n4620, ZN => n4623);
   U2464 : XNOR2_X1 port map( A => n4623, B => n4622, ZN => n4643);
   U2465 : NAND2_X1 port map( A1 => n4625, A2 => n4624, ZN => n4629);
   U2466 : XNOR2_X1 port map( A => n4627, B => n4626, ZN => n4628);
   U2467 : XNOR2_X1 port map( A => n4629, B => n4628, ZN => n4644);
   U2468 : NAND2_X1 port map( A1 => n4643, A2 => n4644, ZN => n4683);
   U2469 : XNOR2_X1 port map( A => n4631, B => n4630, ZN => n4770);
   U2470 : INV_X1 port map( A => n4770, ZN => n4642);
   U2471 : MUX2_X1 port map( A => n4490, B => n8577, S => n395, Z => n4634);
   U2472 : MUX2_X1 port map( A => n4607, B => n8595, S => n2638, Z => n4633);
   U2473 : NAND2_X1 port map( A1 => n4634, A2 => n4633, ZN => n4640);
   U2474 : INV_X1 port map( A => n4640, ZN => n4637);
   U2475 : MUX2_X1 port map( A => n4975, B => n8012, S => n8333, Z => n4636);
   U2476 : MUX2_X1 port map( A => n8455, B => n8553, S => n8564, Z => n4635);
   U2477 : NOR2_X1 port map( A1 => n4636, A2 => n4635, ZN => n4638);
   U2478 : NAND2_X1 port map( A1 => n4637, A2 => n4638, ZN => n4768);
   U2479 : INV_X1 port map( A => n4768, ZN => n4641);
   U2480 : INV_X1 port map( A => n4638, ZN => n4639);
   U2481 : NAND2_X1 port map( A1 => n4640, A2 => n4639, ZN => n4767);
   U2482 : OAI21_X1 port map( B1 => n4642, B2 => n4641, A => n4767, ZN => n4684
                           );
   U2483 : NAND2_X1 port map( A1 => n4683, A2 => n4684, ZN => n4647);
   U2484 : INV_X1 port map( A => n4643, ZN => n4646);
   U2485 : INV_X1 port map( A => n4644, ZN => n4645);
   U2486 : NAND2_X1 port map( A1 => n4646, A2 => n4645, ZN => n4682);
   U2487 : NAND2_X1 port map( A1 => n4647, A2 => n4682, ZN => n4686);
   U2488 : XNOR2_X1 port map( A => n4648, B => n4686, ZN => n4943);
   U2489 : NAND2_X1 port map( A1 => n4650, A2 => n4649, ZN => n4653);
   U2490 : INV_X1 port map( A => n4651, ZN => n4652);
   U2491 : XNOR2_X1 port map( A => n4653, B => n4652, ZN => n4676);
   U2492 : INV_X1 port map( A => n4676, ZN => n4663);
   U2493 : MUX2_X1 port map( A => n8445, B => n6740, S => n8324, Z => n4655);
   U2494 : MUX2_X1 port map( A => n8459, B => n8434, S => n8328, Z => n4654);
   U2495 : NAND2_X1 port map( A1 => n4655, A2 => n4654, ZN => n4752);
   U2496 : MUX2_X1 port map( A => n7946, B => n7947, S => n204, Z => n4657);
   U2497 : NAND2_X1 port map( A1 => n5781, A2 => n8327, ZN => n4656);
   U2498 : NAND2_X1 port map( A1 => n4491, A2 => n8354, ZN => n4749);
   U2499 : NOR2_X1 port map( A1 => n4659, A2 => n4749, ZN => n4661);
   U2500 : INV_X1 port map( A => n4749, ZN => n4660);
   U2501 : OAI22_X1 port map( A1 => n4752, A2 => n4661, B1 => n4660, B2 => 
                           n4750, ZN => n4675);
   U2502 : INV_X1 port map( A => n4675, ZN => n4662);
   U2503 : NAND2_X1 port map( A1 => n4663, A2 => n4662, ZN => n4745);
   U2504 : MUX2_X1 port map( A => n8547, B => n8546, S => n8564, Z => n4665);
   U2505 : INV_X1 port map( A => n8552, ZN => n6103);
   U2506 : MUX2_X1 port map( A => n5878, B => n6102, S => n8401, Z => n4664);
   U2507 : NAND2_X1 port map( A1 => n4665, A2 => n4664, ZN => n4670);
   U2508 : MUX2_X1 port map( A => n8510, B => n4867, S => n6109, Z => n4667);
   U2509 : MUX2_X1 port map( A => n8454, B => n8516, S => n362, Z => n4666);
   U2510 : NAND2_X1 port map( A1 => n4667, A2 => n4666, ZN => n4671);
   U2511 : NAND2_X1 port map( A1 => n4670, A2 => n4671, ZN => n8020);
   U2512 : MUX2_X1 port map( A => n6714, B => n6888, S => n381, Z => n4669);
   U2513 : MUX2_X1 port map( A => n6715, B => n6887, S => n395, Z => n4668);
   U2514 : AND2_X1 port map( A1 => n4669, A2 => n4668, ZN => n8022);
   U2515 : NAND2_X1 port map( A1 => n8020, A2 => n8022, ZN => n4674);
   U2516 : INV_X1 port map( A => n4670, ZN => n4673);
   U2517 : INV_X1 port map( A => n4671, ZN => n4672);
   U2518 : NAND2_X1 port map( A1 => n4673, A2 => n4672, ZN => n8021);
   U2519 : NAND2_X1 port map( A1 => n4674, A2 => n8021, ZN => n4747);
   U2520 : NAND2_X1 port map( A1 => n4745, A2 => n4747, ZN => n4677);
   U2521 : NAND2_X1 port map( A1 => n4676, A2 => n4675, ZN => n4746);
   U2522 : NAND2_X1 port map( A1 => n4679, A2 => n4678, ZN => n4680);
   U2523 : XNOR2_X1 port map( A => n4681, B => n4680, ZN => n4936);
   U2524 : NAND2_X1 port map( A1 => n4683, A2 => n4682, ZN => n4685);
   U2525 : XNOR2_X1 port map( A => n4685, B => n4684, ZN => n4938);
   U2526 : FA_X1 port map( A => n4935, B => n4936, CI => n4938, CO => n4944, S 
                           => n_1129);
   U2527 : NOR2_X1 port map( A1 => n4943, A2 => n4944, ZN => n4949);
   U2528 : NAND2_X1 port map( A1 => n4687, A2 => n4686, ZN => n4688);
   U2529 : AND2_X1 port map( A1 => n4689, A2 => n4688, ZN => n5022);
   U2530 : NAND2_X1 port map( A1 => n4691, A2 => n4690, ZN => n4693);
   U2531 : NAND2_X1 port map( A1 => n4695, A2 => n4694, ZN => n5007);
   U2532 : NAND2_X1 port map( A1 => n5007, A2 => n5006, ZN => n5011);
   U2533 : INV_X1 port map( A => n5011, ZN => n4701);
   U2534 : MUX2_X1 port map( A => n6714, B => n6888, S => n390, Z => n4697);
   U2535 : MUX2_X1 port map( A => n6715, B => n6887, S => n6606, Z => n4696);
   U2536 : MUX2_X1 port map( A => n5898, B => n6249, S => n373, Z => n4699);
   U2537 : MUX2_X1 port map( A => n8454, B => n8516, S => n379, Z => n4698);
   U2538 : NAND2_X1 port map( A1 => n4699, A2 => n4698, ZN => n5005);
   U2539 : XNOR2_X1 port map( A => n5008, B => n5005, ZN => n4700);
   U2540 : XNOR2_X1 port map( A => n4701, B => n4700, ZN => n4715);
   U2541 : MUX2_X1 port map( A => n5845, B => n5844, S => n204, Z => n4703);
   U2542 : MUX2_X1 port map( A => n6103, B => n6102, S => B_SIG_9_port, Z => 
                           n4702);
   U2543 : NAND2_X1 port map( A1 => n4703, A2 => n4702, ZN => n4709);
   U2544 : INV_X1 port map( A => n4709, ZN => n4707);
   U2545 : MUX2_X1 port map( A => n7946, B => n7947, S => n359, Z => n4705);
   U2546 : NAND2_X1 port map( A1 => n5781, A2 => n356, ZN => n4704);
   U2547 : NAND2_X1 port map( A1 => n4705, A2 => n4704, ZN => n4708);
   U2548 : INV_X1 port map( A => n4708, ZN => n4706);
   U2549 : NAND2_X1 port map( A1 => n4707, A2 => n4706, ZN => n5003);
   U2550 : NAND2_X1 port map( A1 => n4709, A2 => n4708, ZN => n5002);
   U2551 : NAND2_X1 port map( A1 => n5003, A2 => n5002, ZN => n4713);
   U2552 : MUX2_X1 port map( A => n4490, B => n8577, S => n8324, Z => n4711);
   U2553 : MUX2_X1 port map( A => n4607, B => n8596, S => n386, Z => n4710);
   U2554 : AND2_X1 port map( A1 => n4711, A2 => n4710, ZN => n5001);
   U2555 : INV_X1 port map( A => n5001, ZN => n4712);
   U2556 : XNOR2_X1 port map( A => n4713, B => n4712, ZN => n4714);
   U2557 : NAND2_X1 port map( A1 => n4715, A2 => n4714, ZN => n4990);
   U2558 : INV_X1 port map( A => n4714, ZN => n4717);
   U2559 : INV_X1 port map( A => n4715, ZN => n4716);
   U2560 : NAND2_X1 port map( A1 => n4717, A2 => n4716, ZN => n4991);
   U2561 : NAND2_X1 port map( A1 => n4990, A2 => n4991, ZN => n5015);
   U2562 : XNOR2_X1 port map( A => n5015, B => n5016, ZN => n4744);
   U2563 : NAND2_X1 port map( A1 => n4718, A2 => n4719, ZN => n4722);
   U2564 : INV_X1 port map( A => n4718, ZN => n4721);
   U2565 : INV_X1 port map( A => n4719, ZN => n4720);
   U2566 : AOI22_X1 port map( A1 => n4723, A2 => n4722, B1 => n4721, B2 => 
                           n4720, ZN => n4734);
   U2568 : XNOR2_X1 port map( A => n4961, B => n8396, ZN => n4724);
   U2569 : NAND2_X1 port map( A1 => n5307, A2 => n4724, ZN => n4726);
   U2570 : INV_X1 port map( A => n4963, ZN => n7010);
   U2571 : NAND2_X1 port map( A1 => n7010, A2 => n395, ZN => n4725);
   U2573 : XNOR2_X2 port map( A => n394, B => n8361, ZN => n5040);
   U2574 : INV_X1 port map( A => n5040, ZN => n6687);
   U2575 : NOR2_X1 port map( A1 => n6687, A2 => n2638, ZN => n4953);
   U2576 : XNOR2_X1 port map( A => n4954, B => n4953, ZN => n4732);
   U2577 : MUX2_X1 port map( A => n8004, B => n8003, S => n8333, Z => n4730);
   U2578 : XNOR2_X1 port map( A => n7945, B => n8002, ZN => n4728);
   U2579 : NAND2_X1 port map( A1 => n4728, A2 => n6264, ZN => n4729);
   U2580 : AND2_X1 port map( A1 => n4730, A2 => n4729, ZN => n4956);
   U2581 : INV_X1 port map( A => n4956, ZN => n4731);
   U2582 : XNOR2_X1 port map( A => n4732, B => n4731, ZN => n4733);
   U2583 : OAI21_X1 port map( B1 => n4423, B2 => n4737, A => n4736, ZN => n4986
                           );
   U2584 : XNOR2_X1 port map( A => n4738, B => n4986, ZN => n5017);
   U2585 : INV_X1 port map( A => n5017, ZN => n4742);
   U2586 : OAI21_X1 port map( B1 => n4741, B2 => n4740, A => n4739, ZN => n5014
                           );
   U2587 : XNOR2_X1 port map( A => n4742, B => n5014, ZN => n4743);
   U2588 : XNOR2_X1 port map( A => n4744, B => n4743, ZN => n5021);
   U2589 : NAND2_X1 port map( A1 => n5022, A2 => n5021, ZN => n4950);
   U2590 : NAND2_X1 port map( A1 => n4746, A2 => n4745, ZN => n4748);
   U2591 : XNOR2_X1 port map( A => n4748, B => n4747, ZN => n4932);
   U2592 : XNOR2_X1 port map( A => n4750, B => n4749, ZN => n4751);
   U2593 : XNOR2_X1 port map( A => n4752, B => n4751, ZN => n4765);
   U2594 : MUX2_X1 port map( A => n8445, B => n6740, S => n386, Z => n4754);
   U2595 : MUX2_X1 port map( A => n8459, B => n8434, S => n8396, Z => n4753);
   U2596 : NAND2_X1 port map( A1 => n4754, A2 => n4753, ZN => n8009);
   U2597 : MUX2_X1 port map( A => n7947, B => n7946, S => B_SIG_9_port, Z => 
                           n4756);
   U2599 : OR2_X1 port map( A1 => n7949, A2 => n7945, ZN => n4755);
   U2600 : NAND2_X1 port map( A1 => n4756, A2 => n4755, ZN => n8010);
   U2601 : NAND2_X1 port map( A1 => n8009, A2 => n8010, ZN => n8008);
   U2602 : NAND2_X1 port map( A1 => n4765, A2 => n8008, ZN => n4766);
   U2603 : OAI21_X1 port map( B1 => n6888, B2 => n8354, A => n6887, ZN => n4761
                           );
   U2604 : MUX2_X1 port map( A => n5398, B => n5397, S => n390, Z => n4762);
   U2605 : NOR2_X1 port map( A1 => n4761, A2 => n4762, ZN => n4757);
   U2606 : MUX2_X1 port map( A => n4867, B => n8535, S => n362, Z => n4760);
   U2607 : NAND2_X1 port map( A1 => n4757, A2 => n4760, ZN => n4774);
   U2608 : MUX2_X1 port map( A => n6714, B => n6888, S => n395, Z => n4759);
   U2609 : MUX2_X1 port map( A => n6715, B => n6887, S => n2638, Z => n4758);
   U2610 : NAND2_X1 port map( A1 => n4759, A2 => n4758, ZN => n4776);
   U2611 : NAND2_X1 port map( A1 => n4774, A2 => n4776, ZN => n4764);
   U2612 : INV_X1 port map( A => n4760, ZN => n4763);
   U2613 : OAI21_X1 port map( B1 => n4763, B2 => n4762, A => n4761, ZN => n4775
                           );
   U2614 : NAND2_X1 port map( A1 => n4764, A2 => n4775, ZN => n8017);
   U2615 : INV_X1 port map( A => n4765, ZN => n8018);
   U2616 : INV_X1 port map( A => n8008, ZN => n8016);
   U2617 : AOI22_X1 port map( A1 => n4766, A2 => n8017, B1 => n8018, B2 => 
                           n8016, ZN => n4934);
   U2618 : NAND2_X1 port map( A1 => n4768, A2 => n4767, ZN => n4769);
   U2619 : XNOR2_X1 port map( A => n4770, B => n4769, ZN => n4931);
   U2620 : XNOR2_X1 port map( A => n4934, B => n4931, ZN => n4771);
   U2621 : XNOR2_X1 port map( A => n4771, B => n4932, ZN => n4926);
   U2622 : NAND2_X1 port map( A1 => n4950, A2 => n4772, ZN => n4773);
   U2623 : NOR2_X1 port map( A1 => n4949, A2 => n4773, ZN => n4942);
   U2624 : NAND2_X1 port map( A1 => n4775, A2 => n4774, ZN => n4777);
   U2625 : XNOR2_X1 port map( A => n4777, B => n4776, ZN => n4802);
   U2626 : MUX2_X1 port map( A => n8488, B => n5395, S => n8564, Z => n4779);
   U2627 : MUX2_X1 port map( A => n5398, B => n5397, S => n376, Z => n4778);
   U2628 : NOR2_X1 port map( A1 => n4779, A2 => n4778, ZN => n4787);
   U2629 : MUX2_X1 port map( A => n8445, B => n6740, S => n395, Z => n4781);
   U2630 : MUX2_X1 port map( A => n8459, B => n8434, S => n8354, Z => n4780);
   U2631 : NAND2_X1 port map( A1 => n4781, A2 => n4780, ZN => n4851);
   U2632 : INV_X1 port map( A => n6740, ZN => n6744);
   U2633 : AOI21_X1 port map( B1 => n6744, B2 => n2638, A => n5033, ZN => n4782
                           );
   U2634 : INV_X1 port map( A => n4782, ZN => n4852);
   U2635 : NAND2_X1 port map( A1 => n4851, A2 => n4852, ZN => n4850);
   U2636 : INV_X1 port map( A => n4787, ZN => n4789);
   U2637 : NAND2_X1 port map( A1 => n4787, A2 => n4782, ZN => n4785);
   U2638 : MUX2_X1 port map( A => n8438, B => n8436, S => n8324, Z => n4784);
   U2639 : MUX2_X1 port map( A => n5878, B => n6102, S => n8328, Z => n4783);
   U2640 : NAND2_X1 port map( A1 => n4784, A2 => n4783, ZN => n4788);
   U2641 : OAI211_X1 port map( C1 => n4851, C2 => n4789, A => n4785, B => n4788
                           , ZN => n4786);
   U2642 : OAI21_X1 port map( B1 => n4787, B2 => n4850, A => n4786, ZN => n4801
                           );
   U2643 : FA_X1 port map( A => n4802, B => n4801, CI => intadd_33_SUM_1_port, 
                           CO => n4927, S => n_1130);
   U2644 : XNOR2_X1 port map( A => n4789, B => n4788, ZN => n4791);
   U2645 : INV_X1 port map( A => n4850, ZN => n4790);
   U2646 : XNOR2_X1 port map( A => n4791, B => n4790, ZN => n4920);
   U2647 : MUX2_X1 port map( A => n4867, B => n8510, S => n6606, Z => n4793);
   U2648 : MUX2_X1 port map( A => n8454, B => n8515, S => n8324, Z => n4792);
   U2649 : NAND2_X1 port map( A1 => n4793, A2 => n4792, ZN => n4860);
   U2650 : INV_X1 port map( A => n4860, ZN => n4800);
   U2651 : MUX2_X1 port map( A => n8547, B => n8546, S => n386, Z => n4795);
   U2652 : MUX2_X1 port map( A => n5878, B => n6102, S => n8396, Z => n4794);
   U2653 : NAND2_X1 port map( A1 => n4795, A2 => n4794, ZN => n4796);
   U2654 : INV_X1 port map( A => n4796, ZN => n4861);
   U2655 : NAND2_X1 port map( A1 => n4796, A2 => n4860, ZN => n4799);
   U2656 : MUX2_X1 port map( A => n7946, B => n7947, S => n362, Z => n4798);
   U2657 : NAND2_X1 port map( A1 => n5781, A2 => n8564, ZN => n4797);
   U2658 : AND2_X1 port map( A1 => n4798, A2 => n4797, ZN => n4858);
   U2659 : AOI22_X1 port map( A1 => n4800, A2 => n4861, B1 => n4799, B2 => 
                           n4858, ZN => n4919);
   U2660 : FA_X1 port map( A => n4920, B => n4919, CI => intadd_33_SUM_0_port, 
                           CO => n4925, S => n_1131);
   U2661 : XNOR2_X1 port map( A => n4802, B => n4801, ZN => n4803);
   U2662 : XNOR2_X1 port map( A => intadd_33_SUM_1_port, B => n4803, ZN => 
                           n4924);
   U2663 : OAI22_X1 port map( A1 => intadd_33_SUM_2_port, A2 => n4927, B1 => 
                           n4925, B2 => n4924, ZN => n4930);
   U2664 : MUX2_X1 port map( A => n5898, B => n8535, S => n386, Z => n4805);
   U2665 : MUX2_X1 port map( A => n8454, B => n8516, S => n381, Z => n4804);
   U2666 : NAND2_X1 port map( A1 => n4805, A2 => n4804, ZN => n4844);
   U2667 : MUX2_X1 port map( A => n7946, B => n7947, S => n376, Z => n4807);
   U2668 : NAND2_X1 port map( A1 => n5781, A2 => n8324, ZN => n4806);
   U2669 : NAND2_X1 port map( A1 => n4807, A2 => n4806, ZN => n4827);
   U2670 : NOR2_X1 port map( A1 => n5846, A2 => n4809, ZN => n6591);
   U2671 : NAND2_X1 port map( A1 => n4810, A2 => n8354, ZN => n4811);
   U2672 : NAND2_X1 port map( A1 => n6591, A2 => n4811, ZN => n4828);
   U2673 : XNOR2_X1 port map( A => n4827, B => n4828, ZN => n4838);
   U2674 : XNOR2_X1 port map( A => n4844, B => n4838, ZN => n4814);
   U2675 : MUX2_X1 port map( A => n8438, B => n8436, S => n395, Z => n4813);
   U2676 : MUX2_X1 port map( A => n5878, B => n6102, S => n8354, Z => n4812);
   U2677 : NAND2_X1 port map( A1 => n4813, A2 => n4812, ZN => n4841);
   U2678 : MUX2_X1 port map( A => n4867, B => n8510, S => n381, Z => n4816);
   U2679 : MUX2_X1 port map( A => n6126, B => n8516, S => n395, Z => n4815);
   U2680 : NAND2_X1 port map( A1 => n4816, A2 => n4815, ZN => n4880);
   U2681 : NOR2_X1 port map( A1 => n6251, A2 => n2638, ZN => n4876);
   U2682 : MUX2_X1 port map( A => n7946, B => n7947, S => n8324, Z => n4819);
   U2683 : NAND2_X1 port map( A1 => n5781, A2 => n386, ZN => n4818);
   U2684 : NAND2_X1 port map( A1 => n4819, A2 => n4818, ZN => n4878);
   U2685 : OAI21_X1 port map( B1 => n4880, B2 => n4876, A => n4878, ZN => n4821
                           );
   U2686 : NAND2_X1 port map( A1 => n4880, A2 => n4876, ZN => n4820);
   U2687 : MUX2_X1 port map( A => n5845, B => n8546, S => n381, Z => n4823);
   U2688 : MUX2_X1 port map( A => n5878, B => n6102, S => n8393, Z => n4822);
   U2689 : NAND2_X1 port map( A1 => n4823, A2 => n4822, ZN => n4855);
   U2690 : MUX2_X1 port map( A => n7946, B => n7947, S => n390, Z => n4825);
   U2691 : NAND2_X1 port map( A1 => n5781, A2 => n376, ZN => n4824);
   U2692 : NAND2_X1 port map( A1 => n4825, A2 => n4824, ZN => n4853);
   U2693 : AND2_X1 port map( A1 => n6264, A2 => n8354, ZN => n4854);
   U2694 : XNOR2_X1 port map( A => n4853, B => n4854, ZN => n4826);
   U2695 : XNOR2_X1 port map( A => n4855, B => n4826, ZN => n4848);
   U2696 : INV_X1 port map( A => n4828, ZN => n4829);
   U2697 : NAND2_X1 port map( A1 => n4827, A2 => n4829, ZN => n4845);
   U2698 : INV_X1 port map( A => n4845, ZN => n4832);
   U2699 : MUX2_X1 port map( A => n4867, B => n8510, S => n8324, Z => n4831);
   U2700 : MUX2_X1 port map( A => n8454, B => n8515, S => n386, Z => n4830);
   U2701 : NAND2_X1 port map( A1 => n4831, A2 => n4830, ZN => n4846);
   U2702 : OAI21_X1 port map( B1 => n4848, B2 => n4832, A => n4846, ZN => n4834
                           );
   U2703 : NAND2_X1 port map( A1 => n4848, A2 => n4832, ZN => n4833);
   U2704 : NAND2_X1 port map( A1 => n4834, A2 => n4833, ZN => n4907);
   U2705 : INV_X1 port map( A => n4907, ZN => n4835);
   U2706 : NAND2_X1 port map( A1 => n4836, A2 => n4835, ZN => n4864);
   U2707 : NAND2_X1 port map( A1 => n4837, A2 => n4898, ZN => n4849);
   U2708 : INV_X1 port map( A => n4841, ZN => n4839);
   U2709 : INV_X1 port map( A => n4838, ZN => n4840);
   U2710 : NAND2_X1 port map( A1 => n4839, A2 => n4840, ZN => n4843);
   U2712 : AOI22_X1 port map( A1 => n4844, A2 => n4843, B1 => n4838, B2 => 
                           n4841, ZN => n4903);
   U2713 : XNOR2_X1 port map( A => n4846, B => n4845, ZN => n4847);
   U2714 : XNOR2_X1 port map( A => n4848, B => n4847, ZN => n4904);
   U2715 : OAI21_X1 port map( B1 => n4852, B2 => n4851, A => n4850, ZN => n4913
                           );
   U2716 : OAI21_X1 port map( B1 => n4855, B2 => n4854, A => n4853, ZN => n4857
                           );
   U2717 : NAND2_X1 port map( A1 => n4855, A2 => n4854, ZN => n4856);
   U2718 : NAND2_X1 port map( A1 => n4857, A2 => n4856, ZN => n4915);
   U2719 : XNOR2_X1 port map( A => n4913, B => n4915, ZN => n4863);
   U2720 : INV_X1 port map( A => n4858, ZN => n4859);
   U2721 : XNOR2_X1 port map( A => n4860, B => n4859, ZN => n4862);
   U2722 : XNOR2_X1 port map( A => n4862, B => n4861, ZN => n4912);
   U2723 : XNOR2_X1 port map( A => n4863, B => n4912, ZN => n4908);
   U2724 : OAI21_X1 port map( B1 => n4864, B2 => n4866, A => n4908, ZN => n4911
                           );
   U2725 : OAI21_X1 port map( B1 => n4866, B2 => n4865, A => n4907, ZN => n4910
                           );
   U2726 : MUX2_X1 port map( A => n4867, B => n8510, S => n395, Z => n4890);
   U2727 : MUX2_X1 port map( A => n6126, B => n8515, S => n2638, Z => n4868);
   U2728 : NAND2_X1 port map( A1 => n4890, A2 => n4868, ZN => n4873);
   U2729 : INV_X1 port map( A => n4873, ZN => n4871);
   U2730 : MUX2_X1 port map( A => n7946, B => n7947, S => n386, Z => n4870);
   U2731 : NAND2_X1 port map( A1 => n5781, A2 => n381, ZN => n4869);
   U2732 : NAND2_X1 port map( A1 => n4870, A2 => n4869, ZN => n4872);
   U2733 : INV_X1 port map( A => n4872, ZN => n4889);
   U2734 : NAND2_X1 port map( A1 => n4871, A2 => n4889, ZN => n4896);
   U2735 : INV_X1 port map( A => n4896, ZN => n4875);
   U2736 : AOI21_X1 port map( B1 => n5395, B2 => n2638, A => n5397, ZN => n4874
                           );
   U2737 : NAND2_X1 port map( A1 => n4873, A2 => n4872, ZN => n4883);
   U2738 : OAI21_X1 port map( B1 => n4875, B2 => n4874, A => n4883, ZN => n4882
                           );
   U2739 : INV_X1 port map( A => n4876, ZN => n4877);
   U2740 : XNOR2_X1 port map( A => n4878, B => n4877, ZN => n4879);
   U2741 : XNOR2_X1 port map( A => n4880, B => n4879, ZN => n4884);
   U2742 : INV_X1 port map( A => n4884, ZN => n4881);
   U2743 : NAND2_X1 port map( A1 => n4882, A2 => n4881, ZN => n4902);
   U2744 : NAND2_X1 port map( A1 => n4884, A2 => n4883, ZN => n4897);
   U2745 : MUX2_X1 port map( A => n7946, B => n7947, S => n381, Z => n4887);
   U2746 : NAND2_X1 port map( A1 => n5781, A2 => n395, ZN => n4886);
   U2747 : AOI21_X1 port map( B1 => n4887, B2 => n4886, A => n5055, ZN => n4888
                           );
   U2748 : OAI21_X1 port map( B1 => n4890, B2 => n4889, A => n4888, ZN => n4891
                           );
   U2749 : NAND2_X1 port map( A1 => n4891, A2 => n8354, ZN => n4895);
   U2750 : NAND2_X1 port map( A1 => n395, A2 => n381, ZN => n4893);
   U2751 : OAI21_X1 port map( B1 => n4893, B2 => n6259, A => n2638, ZN => n4894
                           );
   U2752 : NAND4_X1 port map( A1 => n4897, A2 => n4896, A3 => n4895, A4 => 
                           n4894, ZN => n4901);
   U2753 : INV_X1 port map( A => n4898, ZN => n4899);
   U2754 : AOI22_X1 port map( A1 => n4902, A2 => n4901, B1 => n4900, B2 => 
                           n4899, ZN => n4906);
   U2755 : NAND2_X1 port map( A1 => n4904, A2 => n4903, ZN => n4905);
   U2756 : OAI211_X1 port map( C1 => n4908, C2 => n4907, A => n4906, B => n4905
                           , ZN => n4909);
   U2757 : INV_X1 port map( A => n4912, ZN => n4916);
   U2758 : INV_X1 port map( A => n4913, ZN => n4914);
   U2759 : OAI21_X1 port map( B1 => n4916, B2 => n4915, A => n4914, ZN => n4918
                           );
   U2760 : NAND2_X1 port map( A1 => n4916, A2 => n4915, ZN => n4917);
   U2761 : NAND2_X1 port map( A1 => n4918, A2 => n4917, ZN => n4923);
   U2762 : XNOR2_X1 port map( A => intadd_33_SUM_0_port, B => n4919, ZN => 
                           n4921);
   U2763 : XNOR2_X1 port map( A => n4921, B => n4920, ZN => n4922);
   U2764 : AOI22_X1 port map( A1 => intadd_33_SUM_2_port, A2 => n4927, B1 => 
                           intadd_33_n1, B2 => n4926, ZN => n4928);
   U2765 : OAI21_X1 port map( B1 => n4930, B2 => n4929, A => n4928, ZN => n4941
                           );
   U2766 : INV_X1 port map( A => n4931, ZN => n4933);
   U2767 : FA_X1 port map( A => n4934, B => n4933, CI => n4932, CO => n4946, S 
                           => n_1132);
   U2768 : INV_X1 port map( A => n4935, ZN => n4937);
   U2769 : XNOR2_X1 port map( A => n4937, B => n4936, ZN => n4939);
   U2770 : XNOR2_X1 port map( A => n4939, B => n4938, ZN => n4945);
   U2771 : NAND2_X1 port map( A1 => n4946, A2 => n4945, ZN => n4940);
   U2772 : NAND3_X1 port map( A1 => n4942, A2 => n4941, A3 => n4940, ZN => 
                           n5029);
   U2773 : INV_X1 port map( A => n4943, ZN => n4948);
   U2774 : INV_X1 port map( A => n4944, ZN => n4947);
   U2775 : OAI22_X1 port map( A1 => n4948, A2 => n4947, B1 => n4945, B2 => 
                           n4946, ZN => n4952);
   U2776 : INV_X1 port map( A => n4949, ZN => n4951);
   U2777 : NAND3_X1 port map( A1 => n4952, A2 => n4951, A3 => n4950, ZN => 
                           n5028);
   U2778 : NAND2_X1 port map( A1 => n4954, A2 => n4953, ZN => n4957);
   U2779 : NOR2_X1 port map( A1 => n4954, A2 => n4953, ZN => n4955);
   U2780 : MUX2_X1 port map( A => n6714, B => n6888, S => n362, Z => n4959);
   U2781 : MUX2_X1 port map( A => n6715, B => n6887, S => n390, Z => n4958);
   U2782 : AND2_X1 port map( A1 => n4959, A2 => n4958, ZN => n5120);
   U2783 : XNOR2_X1 port map( A => n5116, B => n4960, ZN => n4972);
   U2784 : NAND2_X1 port map( A1 => n4962, A2 => n4961, ZN => n5030);
   U2785 : MUX2_X1 port map( A => n8593, B => n7122, S => n381, Z => n4964);
   U2786 : NAND2_X1 port map( A1 => n4965, A2 => n4964, ZN => n5104);
   U2787 : NAND2_X1 port map( A1 => n8003, A2 => n6109, ZN => n4967);
   U2788 : NAND2_X1 port map( A1 => n8004, A2 => n8362, ZN => n4966);
   U2789 : NAND2_X1 port map( A1 => n4967, A2 => n4966, ZN => n4970);
   U2790 : XNOR2_X1 port map( A => B_SIG_9_port, B => n8002, ZN => n4968);
   U2791 : NAND2_X1 port map( A1 => n6264, A2 => n4968, ZN => n4969);
   U2792 : NAND2_X1 port map( A1 => n4970, A2 => n4969, ZN => n5103);
   U2793 : INV_X1 port map( A => n5103, ZN => n4971);
   U2794 : XNOR2_X1 port map( A => n5104, B => n4971, ZN => n5117);
   U2795 : XNOR2_X1 port map( A => n4972, B => n5117, ZN => n4985);
   U2796 : MUX2_X1 port map( A => n8488, B => n5395, S => n356, Z => n4974);
   U2797 : MUX2_X1 port map( A => n5398, B => n5397, S => n373, Z => n4973);
   U2798 : NOR2_X1 port map( A1 => n4974, A2 => n4973, ZN => n4978);
   U2799 : MUX2_X1 port map( A => n4975, B => n8012, S => n8392, Z => n4977);
   U2800 : MUX2_X1 port map( A => n5794, B => n8553, S => n204, Z => n4976);
   U2801 : NOR2_X1 port map( A1 => n4977, A2 => n4976, ZN => n4979);
   U2802 : NAND2_X1 port map( A1 => n4978, A2 => n4979, ZN => n5114);
   U2803 : NAND2_X1 port map( A1 => n5114, A2 => n5112, ZN => n4983);
   U2804 : MUX2_X1 port map( A => n4490, B => n8577, S => n6606, Z => n4981);
   U2805 : MUX2_X1 port map( A => n4607, B => n8596, S => n8324, Z => n4980);
   U2806 : AND2_X1 port map( A1 => n4981, A2 => n4980, ZN => n5111);
   U2807 : INV_X1 port map( A => n5111, ZN => n4982);
   U2808 : XNOR2_X1 port map( A => n4983, B => n4982, ZN => n4984);
   U2809 : NAND2_X1 port map( A1 => n4985, A2 => n4984, ZN => n5159);
   U2810 : NAND2_X1 port map( A1 => n5160, A2 => n5159, ZN => n4989);
   U2811 : NAND2_X1 port map( A1 => n4988, A2 => n4987, ZN => n5158);
   U2812 : XNOR2_X1 port map( A => n4989, B => n5158, ZN => n5171);
   U2813 : NAND2_X1 port map( A1 => n5014, A2 => n4990, ZN => n4992);
   U2814 : NAND2_X1 port map( A1 => n4992, A2 => n4991, ZN => n5172);
   U2815 : NAND2_X2 port map( A1 => n5040, A2 => n8369, ZN => n7080);
   U2816 : INV_X1 port map( A => n7080, ZN => n7215);
   U2817 : NAND2_X1 port map( A1 => n7215, A2 => n2638, ZN => n5101);
   U2819 : NAND2_X1 port map( A1 => n5101, A2 => n7324, ZN => n4995);
   U2820 : XNOR2_X1 port map( A => n377, B => n4892, ZN => n4994);
   U2821 : OAI22_X1 port map( A1 => mult_x_19_n4, A2 => n4994, B1 => n7949, B2 
                           => n8394, ZN => n5095);
   U2822 : INV_X1 port map( A => n5095, ZN => n5102);
   U2824 : BUF_X2 port map( A => n384, Z => n6229);
   U2825 : NAND2_X2 port map( A1 => n5040, A2 => n6229, ZN => n7195);
   U2826 : MUX2_X1 port map( A => n7195, B => n7080, S => n395, Z => n5099);
   U2827 : NOR2_X1 port map( A1 => n394, A2 => n358, ZN => n4997);
   U2829 : MUX2_X1 port map( A => n7324, B => n8465, S => n8354, Z => n4998);
   U2830 : NAND2_X1 port map( A1 => n5099, A2 => n4998, ZN => n4999);
   U2831 : INV_X1 port map( A => n5126, ZN => n5128);
   U2832 : NAND2_X1 port map( A1 => n5002, A2 => n5001, ZN => n5004);
   U2833 : NAND2_X1 port map( A1 => n5004, A2 => n5003, ZN => n5127);
   U2834 : XNOR2_X1 port map( A => n5128, B => n5127, ZN => n5013);
   U2835 : INV_X1 port map( A => n5005, ZN => n5012);
   U2836 : NAND3_X1 port map( A1 => n5007, A2 => n5006, A3 => n5005, ZN => 
                           n5010);
   U2837 : AOI22_X1 port map( A1 => n5012, A2 => n5011, B1 => n5010, B2 => 
                           n5009, ZN => n5131);
   U2838 : XNOR2_X1 port map( A => n5013, B => n5131, ZN => n5173);
   U2839 : INV_X1 port map( A => n5174, ZN => n5026);
   U2840 : XNOR2_X1 port map( A => n5015, B => n5014, ZN => n5020);
   U2841 : INV_X1 port map( A => n5175, ZN => n5025);
   U2842 : INV_X1 port map( A => n5021, ZN => n5024);
   U2843 : INV_X1 port map( A => n5022, ZN => n5023);
   U2844 : AOI22_X1 port map( A1 => n5026, A2 => n5025, B1 => n5024, B2 => 
                           n5023, ZN => n5027);
   U2845 : NAND3_X1 port map( A1 => n5029, A2 => n5028, A3 => n5027, ZN => 
                           n7927);
   U2847 : INV_X1 port map( A => n6811, ZN => n7012);
   U2848 : NAND2_X1 port map( A1 => n4360, A2 => n8324, ZN => n5083);
   U2849 : OAI21_X1 port map( B1 => n8530, B2 => n8324, A => n5083, ZN => n5037
                           );
   U2850 : NAND2_X1 port map( A1 => n7123, A2 => n8328, ZN => n5032);
   U2851 : NAND2_X1 port map( A1 => n6812, A2 => n386, ZN => n5031);
   U2852 : NAND2_X1 port map( A1 => n5032, A2 => n5031, ZN => n5085);
   U2853 : NAND2_X1 port map( A1 => n5037, A2 => n8441, ZN => n5035);
   U2854 : BUF_X2 port map( A => n5142, Z => n6702);
   U2855 : AND2_X1 port map( A1 => n6702, A2 => n8354, ZN => n5036);
   U2856 : MUX2_X1 port map( A => n5034, B => n5033, S => n8327, Z => n5090);
   U2857 : AOI21_X1 port map( B1 => n5035, B2 => n5036, A => n5090, ZN => n5039
                           );
   U2858 : MUX2_X1 port map( A => n8445, B => n6740, S => n204, Z => n5091);
   U2859 : INV_X1 port map( A => n5036, ZN => n5088);
   U2860 : AND3_X1 port map( A1 => n5085, A2 => n5037, A3 => n5088, ZN => n5038
                           );
   U2861 : AOI21_X1 port map( B1 => n5039, B2 => n5091, A => n5038, ZN => n5185
                           );
   U2863 : XNOR2_X1 port map( A => n8396, B => n6229, ZN => n5042);
   U2864 : NAND2_X1 port map( A1 => n5041, A2 => n5042, ZN => n5043);
   U2865 : MUX2_X1 port map( A => n7946, B => n7947, S => n360, Z => n5045);
   U2866 : NAND2_X1 port map( A1 => n5781, A2 => n377, ZN => n5044);
   U2867 : NAND2_X1 port map( A1 => n5045, A2 => n5044, ZN => n5046);
   U2868 : NAND2_X1 port map( A1 => n5047, A2 => n5046, ZN => n5077);
   U2869 : MUX2_X1 port map( A => n4607, B => n8596, S => n376, Z => n5079);
   U2870 : AND2_X1 port map( A1 => n5077, A2 => n5079, ZN => n5048);
   U2871 : MUX2_X1 port map( A => n4490, B => n8577, S => n8564, Z => n5080);
   U2872 : NOR2_X1 port map( A1 => n5047, A2 => n5046, ZN => n5076);
   U2873 : AOI21_X1 port map( B1 => n5048, B2 => n5080, A => n5076, ZN => n5184
                           );
   U2874 : XNOR2_X1 port map( A => n5185, B => n5184, ZN => n5061);
   U2875 : MUX2_X1 port map( A => n8438, B => n8436, S => n373, Z => n5050);
   U2876 : MUX2_X1 port map( A => n5878, B => n6102, S => n8392, Z => n5049);
   U2877 : NAND2_X1 port map( A1 => n5050, A2 => n5049, ZN => n5074);
   U2878 : MUX2_X1 port map( A => n6715, B => n6243, S => n362, Z => n5054);
   U2879 : XNOR2_X1 port map( A => n7945, B => n6244, ZN => n5052);
   U2880 : NAND2_X1 port map( A1 => n5052, A2 => n7861, ZN => n5053);
   U2881 : NAND2_X1 port map( A1 => n5054, A2 => n5053, ZN => n5073);
   U2882 : MUX2_X1 port map( A => n6126, B => n8516, S => n356, Z => n5058);
   U2883 : INV_X1 port map( A => n5055, ZN => n5835);
   U2884 : XNOR2_X1 port map( A => n8394, B => n5848, ZN => n5056);
   U2885 : NAND2_X1 port map( A1 => n5835, A2 => n5056, ZN => n5057);
   U2886 : NAND2_X1 port map( A1 => n5058, A2 => n5057, ZN => n5072);
   U2887 : AOI21_X1 port map( B1 => n5074, B2 => n5073, A => n5072, ZN => n5060
                           );
   U2888 : NOR2_X1 port map( A1 => n5074, A2 => n5073, ZN => n5059);
   U2889 : NOR2_X1 port map( A1 => n5060, A2 => n5059, ZN => n5186);
   U2890 : XNOR2_X1 port map( A => n5061, B => n5186, ZN => n5183);
   U2891 : MUX2_X1 port map( A => n4487, B => n7325, S => n386, Z => n5063);
   U2892 : MUX2_X1 port map( A => n7324, B => n8465, S => n8396, Z => n5062);
   U2893 : NAND2_X1 port map( A1 => n5063, A2 => n5062, ZN => n5187);
   U2894 : INV_X1 port map( A => n5187, ZN => n5066);
   U2895 : MUX2_X1 port map( A => n8438, B => n8436, S => n356, Z => n5065);
   U2896 : MUX2_X1 port map( A => n5878, B => n6102, S => n4381, Z => n5064);
   U2897 : NAND2_X1 port map( A1 => n5065, A2 => n5064, ZN => n5188);
   U2898 : XNOR2_X1 port map( A => n5066, B => n5188, ZN => n5071);
   U2899 : MUX2_X1 port map( A => n7123, B => n7122, S => n8324, Z => n5067);
   U2900 : NAND2_X1 port map( A1 => n5068, A2 => n5067, ZN => n5352);
   U2901 : MUX2_X1 port map( A => n8445, B => n6740, S => n379, Z => n5070);
   U2902 : MUX2_X1 port map( A => n8459, B => n8434, S => n8351, Z => n5069);
   U2903 : NAND2_X1 port map( A1 => n5070, A2 => n5069, ZN => n5353);
   U2904 : NAND2_X1 port map( A1 => n5353, A2 => n5352, ZN => n5211);
   U2905 : OAI21_X1 port map( B1 => n5352, B2 => n5353, A => n5211, ZN => n5202
                           );
   U2907 : XNOR2_X1 port map( A => n5073, B => n5072, ZN => n5075);
   U2908 : XNOR2_X1 port map( A => n5075, B => n5074, ZN => n5164);
   U2909 : INV_X1 port map( A => n5076, ZN => n5078);
   U2910 : NAND2_X1 port map( A1 => n5078, A2 => n5077, ZN => n5082);
   U2911 : NAND2_X1 port map( A1 => n5080, A2 => n5079, ZN => n5081);
   U2912 : XNOR2_X1 port map( A => n5082, B => n5081, ZN => n5163);
   U2913 : NAND3_X1 port map( A1 => n5085, A2 => n8479, A3 => n8350, ZN => 
                           n5087);
   U2914 : INV_X1 port map( A => n5083, ZN => n5084);
   U2915 : NAND2_X1 port map( A1 => n8441, A2 => n5084, ZN => n5086);
   U2916 : NAND2_X1 port map( A1 => n5087, A2 => n5086, ZN => n5089);
   U2917 : XNOR2_X1 port map( A => n5089, B => n5088, ZN => n5094);
   U2918 : INV_X1 port map( A => n5090, ZN => n5092);
   U2919 : NAND2_X1 port map( A1 => n5092, A2 => n5091, ZN => n5093);
   U2920 : XNOR2_X1 port map( A => n5094, B => n5093, ZN => n5162);
   U2921 : NAND2_X1 port map( A1 => n7324, A2 => n8354, ZN => n5096);
   U2922 : AND2_X1 port map( A1 => n5096, A2 => n5095, ZN => n5098);
   U2923 : NAND2_X1 port map( A1 => n7080, A2 => n7324, ZN => n7444);
   U2924 : OAI22_X1 port map( A1 => n2638, A2 => n8465, B1 => n7324, B2 => 
                           n8354, ZN => n5097);
   U2925 : AOI21_X1 port map( B1 => n5098, B2 => n7444, A => n5097, ZN => n5100
                           );
   U2926 : NAND2_X1 port map( A1 => n5100, A2 => n5099, ZN => n5106);
   U2927 : NAND3_X1 port map( A1 => n5102, A2 => n5101, A3 => n7324, ZN => 
                           n5107);
   U2928 : AND2_X1 port map( A1 => n5107, A2 => n5106, ZN => n5105);
   U2929 : NAND2_X1 port map( A1 => n5105, A2 => n5108, ZN => n5148);
   U2930 : INV_X1 port map( A => n5106, ZN => n5110);
   U2931 : INV_X1 port map( A => n5107, ZN => n5109);
   U2932 : OAI21_X1 port map( B1 => n5110, B2 => n5109, A => n4472, ZN => n5149
                           );
   U2933 : NAND2_X1 port map( A1 => n5148, A2 => n5149, ZN => n5115);
   U2934 : NAND2_X1 port map( A1 => n5112, A2 => n5111, ZN => n5113);
   U2935 : XNOR2_X1 port map( A => n5115, B => n4405, ZN => n5125);
   U2937 : NAND2_X1 port map( A1 => n5117, A2 => n4499, ZN => n5121);
   U2938 : INV_X1 port map( A => n5117, ZN => n5119);
   U2939 : INV_X1 port map( A => n4499, ZN => n5118);
   U2940 : AOI22_X1 port map( A1 => n5121, A2 => n5120, B1 => n5119, B2 => 
                           n5118, ZN => n5124);
   U2941 : INV_X1 port map( A => n5124, ZN => n5122);
   U2942 : NAND2_X1 port map( A1 => n8453, A2 => n5122, ZN => n5155);
   U2943 : NAND2_X1 port map( A1 => n5124, A2 => n5125, ZN => n5154);
   U2944 : NAND2_X1 port map( A1 => n5126, A2 => n5127, ZN => n5130);
   U2945 : INV_X1 port map( A => n5127, ZN => n5129);
   U2947 : NAND2_X1 port map( A1 => n5154, A2 => n5156, ZN => n5132);
   U2948 : AND2_X1 port map( A1 => n5155, A2 => n5132, ZN => n5264);
   U2949 : MUX2_X1 port map( A => n6888, B => n6714, S => B_SIG_9_port, Z => 
                           n5134);
   U2950 : MUX2_X1 port map( A => n6887, B => n6715, S => n6109, Z => n5133);
   U2951 : NAND2_X1 port map( A1 => n5134, A2 => n5133, ZN => n5238);
   U2952 : MUX2_X1 port map( A => n5898, B => n6249, S => n377, Z => n5136);
   U2953 : MUX2_X1 port map( A => n8454, B => n8515, S => n359, Z => n5135);
   U2954 : NAND2_X1 port map( A1 => n5136, A2 => n5135, ZN => n5240);
   U2955 : XNOR2_X1 port map( A => n5238, B => n5240, ZN => n5139);
   U2956 : MUX2_X1 port map( A => n4490, B => n8577, S => n362, Z => n5138);
   U2957 : MUX2_X1 port map( A => n4607, B => n8595, S => n390, Z => n5137);
   U2958 : AND2_X1 port map( A1 => n5138, A2 => n5137, ZN => n5242);
   U2959 : XNOR2_X1 port map( A => n5139, B => n5242, ZN => n5146);
   U2960 : NAND2_X2 port map( A1 => n5142, A2 => n8353, ZN => n7053);
   U2961 : OAI21_X1 port map( B1 => n7053, B2 => n8354, A => n4462, ZN => n5216
                           );
   U2962 : MUX2_X1 port map( A => n7946, B => n7947, S => n372, Z => n5141);
   U2963 : NAND2_X1 port map( A1 => n5781, A2 => n360, ZN => n5140);
   U2964 : NAND2_X1 port map( A1 => n5141, A2 => n5140, ZN => n5213);
   U2965 : INV_X1 port map( A => n5213, ZN => n5217);
   U2966 : XNOR2_X1 port map( A => n5216, B => n5217, ZN => n5145);
   U2967 : BUF_X2 port map( A => n5273, Z => n6705);
   U2968 : MUX2_X1 port map( A => n8501, B => n7053, S => n395, Z => n5214);
   U2971 : NAND2_X2 port map( A1 => n6227, A2 => n6706, ZN => n7054);
   U2972 : BUF_X2 port map( A => n7054, Z => n7198);
   U2973 : MUX2_X1 port map( A => n4462, B => n7198, S => n8354, Z => n5143);
   U2974 : NAND2_X1 port map( A1 => n5214, A2 => n5143, ZN => n5144);
   U2975 : XNOR2_X1 port map( A => n5145, B => n5144, ZN => n5147);
   U2976 : NAND2_X1 port map( A1 => n5146, A2 => n5147, ZN => n5207);
   U2977 : NAND2_X1 port map( A1 => n5207, A2 => n5205, ZN => n5152);
   U2978 : XNOR2_X1 port map( A => n5152, B => n5151, ZN => n5178);
   U2980 : XNOR2_X1 port map( A => n4407, B => n5156, ZN => n5169);
   U2981 : NAND2_X1 port map( A1 => n5159, A2 => n5158, ZN => n5161);
   U2982 : FA_X1 port map( A => n5164, B => n5163, CI => n5162, CO => n5181, S 
                           => n5167);
   U2983 : OAI21_X1 port map( B1 => n4409, B2 => n4477, A => n5167, ZN => n5166
                           );
   U2984 : NAND2_X1 port map( A1 => n4409, A2 => n4477, ZN => n5165);
   U2985 : XNOR2_X1 port map( A => n5168, B => n5167, ZN => n5170);
   U2986 : XNOR2_X1 port map( A => n5169, B => n5170, ZN => n5251);
   U2987 : AOI22_X1 port map( A1 => n5251, A2 => n5252, B1 => n5174, B2 => 
                           n5175, ZN => n5249);
   U2988 : INV_X1 port map( A => n5264, ZN => n5176);
   U2989 : NAND2_X1 port map( A1 => n5177, A2 => n5176, ZN => n5180);
   U2990 : OR2_X1 port map( A1 => n5179, A2 => n5178, ZN => n5262);
   U2991 : NAND2_X1 port map( A1 => n5180, A2 => n5262, ZN => n5266);
   U2992 : FA_X1 port map( A => n5186, B => n5185, CI => n5184, CO => n5369, S 
                           => n_1133);
   U2993 : NAND2_X1 port map( A1 => n5188, A2 => n5187, ZN => n5200);
   U2994 : NOR2_X1 port map( A1 => n5188, A2 => n5187, ZN => n5203);
   U2995 : AOI21_X1 port map( B1 => n5202, B2 => n5200, A => n5203, ZN => n5198
                           );
   U2996 : MUX2_X1 port map( A => n6715, B => n6887, S => n8327, Z => n5191);
   U2997 : XNOR2_X1 port map( A => n8351, B => n6244, ZN => n5189);
   U2998 : NAND2_X1 port map( A1 => n7861, A2 => n5189, ZN => n5190);
   U2999 : NAND2_X1 port map( A1 => n5191, A2 => n5190, ZN => n5281);
   U3000 : MUX2_X1 port map( A => n8454, B => n8515, S => n377, Z => n5194);
   U3001 : XNOR2_X1 port map( A => n8356, B => n360, ZN => n5192);
   U3002 : NAND2_X1 port map( A1 => n5835, A2 => n5192, ZN => n5193);
   U3003 : NAND2_X1 port map( A1 => n5194, A2 => n5193, ZN => n5280);
   U3004 : XNOR2_X1 port map( A => n5281, B => n5280, ZN => n5197);
   U3005 : MUX2_X1 port map( A => n8577, B => n4490, S => n6109, Z => n5196);
   U3006 : MUX2_X1 port map( A => n4607, B => n8596, S => n362, Z => n5195);
   U3007 : NAND2_X1 port map( A1 => n5196, A2 => n5195, ZN => n5282);
   U3008 : XNOR2_X1 port map( A => n5197, B => n5282, ZN => n5199);
   U3009 : NAND2_X1 port map( A1 => n5198, A2 => n5199, ZN => n5366);
   U3010 : INV_X1 port map( A => n5199, ZN => n5201);
   U3011 : OAI211_X1 port map( C1 => n5203, C2 => n5202, A => n5201, B => n5200
                           , ZN => n5367);
   U3012 : NAND2_X1 port map( A1 => n5366, A2 => n5367, ZN => n5204);
   U3013 : XNOR2_X1 port map( A => n5369, B => n5204, ZN => n5376);
   U3014 : XNOR2_X1 port map( A => n5376, B => n5374, ZN => n5247);
   U3015 : NAND2_X1 port map( A1 => n5206, A2 => n5205, ZN => n5208);
   U3016 : NAND2_X1 port map( A1 => n5208, A2 => n5207, ZN => n5335);
   U3017 : MUX2_X1 port map( A => n8438, B => n8436, S => n359, Z => n5210);
   U3018 : MUX2_X1 port map( A => n5878, B => n6102, S => n8326, Z => n5209);
   U3019 : NAND2_X1 port map( A1 => n5210, A2 => n5209, ZN => n5351);
   U3020 : XNOR2_X1 port map( A => n5211, B => n5351, ZN => n5220);
   U3021 : OAI22_X1 port map( A1 => n2638, A2 => n7198, B1 => n4462, B2 => 
                           n8354, ZN => n5212);
   U3022 : AOI21_X1 port map( B1 => n5216, B2 => n5213, A => n5212, ZN => n5215
                           );
   U3023 : NAND2_X1 port map( A1 => n5215, A2 => n5214, ZN => n5349);
   U3024 : INV_X1 port map( A => n5216, ZN => n5218);
   U3025 : NAND2_X1 port map( A1 => n5218, A2 => n5217, ZN => n5348);
   U3026 : NAND2_X1 port map( A1 => n5349, A2 => n5348, ZN => n5219);
   U3027 : XNOR2_X1 port map( A => n5220, B => n5219, ZN => n5334);
   U3028 : XNOR2_X1 port map( A => n5335, B => n5334, ZN => n5246);
   U3029 : MUX2_X1 port map( A => n4461, B => n7054, S => n8393, Z => n5223);
   U3030 : XNOR2_X1 port map( A => n8396, B => n4401, ZN => n5221);
   U3031 : NAND2_X1 port map( A1 => n6702, A2 => n5221, ZN => n5222);
   U3032 : NAND2_X1 port map( A1 => n5223, A2 => n5222, ZN => n5296);
   U3033 : MUX2_X1 port map( A => n7946, B => n7947, S => n363, Z => n5225);
   U3034 : NAND2_X1 port map( A1 => n5781, A2 => n372, ZN => n5224);
   U3035 : NAND2_X1 port map( A1 => n5225, A2 => n5224, ZN => n5297);
   U3036 : XNOR2_X1 port map( A => n5296, B => n5297, ZN => n5229);
   U3037 : INV_X1 port map( A => n7195, ZN => n7216);
   U3038 : MUX2_X1 port map( A => n7216, B => n7215, S => n8324, Z => n5228);
   U3039 : INV_X1 port map( A => n6688, ZN => n6460);
   U3040 : MUX2_X1 port map( A => n6460, B => n5226, S => n386, Z => n5227);
   U3041 : NOR2_X1 port map( A1 => n5228, A2 => n5227, ZN => n5295);
   U3042 : XNOR2_X1 port map( A => n5229, B => n5295, ZN => n5234);
   U3043 : MUX2_X1 port map( A => n8445, B => n6740, S => n373, Z => n5321);
   U3044 : MUX2_X1 port map( A => n8459, B => n8434, S => n8392, Z => n5320);
   U3045 : NAND2_X1 port map( A1 => n5321, A2 => n5320, ZN => n5233);
   U3046 : MUX2_X1 port map( A => n8593, B => n7122, S => n6606, Z => n5231);
   U3047 : XNOR2_X1 port map( A => n8403, B => n390, ZN => n5230);
   U3048 : NAND2_X1 port map( A1 => n5307, A2 => n5230, ZN => n5315);
   U3049 : NAND2_X1 port map( A1 => n5231, A2 => n5315, ZN => n5323);
   U3050 : XNOR2_X1 port map( A => n8359, B => n383, ZN => n5508);
   U3051 : NAND2_X1 port map( A1 => n6595, A2 => n8354, ZN => n5324);
   U3052 : XNOR2_X1 port map( A => n5323, B => n5324, ZN => n5232);
   U3053 : XNOR2_X1 port map( A => n5233, B => n5232, ZN => n5235);
   U3054 : NAND2_X1 port map( A1 => n5234, A2 => n5235, ZN => n5363);
   U3055 : INV_X1 port map( A => n5234, ZN => n5237);
   U3057 : NAND2_X1 port map( A1 => n5237, A2 => n8430, ZN => n5362);
   U3058 : NAND2_X1 port map( A1 => n5363, A2 => n5362, ZN => n5245);
   U3059 : INV_X1 port map( A => n5238, ZN => n5244);
   U3060 : INV_X1 port map( A => n5242, ZN => n5239);
   U3061 : NAND2_X1 port map( A1 => n5239, A2 => n5240, ZN => n5243);
   U3062 : INV_X1 port map( A => n5240, ZN => n5241);
   U3063 : AOI22_X1 port map( A1 => n5244, A2 => n5243, B1 => n5242, B2 => 
                           n5241, ZN => n5360);
   U3064 : XNOR2_X1 port map( A => n5245, B => n5360, ZN => n5333);
   U3066 : XNOR2_X1 port map( A => n5247, B => n4457, ZN => n5259);
   U3067 : NAND2_X1 port map( A1 => n5266, A2 => n5259, ZN => n5248);
   U3068 : OAI211_X1 port map( C1 => n5265, C2 => n5253, A => n5249, B => n5248
                           , ZN => n7929);
   U3069 : INV_X1 port map( A => n7929, ZN => n5250);
   U3070 : NAND2_X1 port map( A1 => n7927, A2 => n5250, ZN => n5380);
   U3071 : INV_X1 port map( A => n5263, ZN => n5258);
   U3072 : INV_X1 port map( A => n5265, ZN => n5257);
   U3073 : INV_X1 port map( A => n5251, ZN => n5255);
   U3074 : INV_X1 port map( A => n5252, ZN => n5254);
   U3075 : NAND3_X1 port map( A1 => n5255, A2 => n5254, A3 => n5253, ZN => 
                           n5267);
   U3076 : AND2_X1 port map( A1 => n5266, A2 => n5267, ZN => n5256);
   U3077 : OAI21_X1 port map( B1 => n5258, B2 => n5257, A => n5256, ZN => n5261
                           );
   U3078 : INV_X1 port map( A => n5259, ZN => n5260);
   U3079 : NAND2_X1 port map( A1 => n5261, A2 => n5260, ZN => n7922);
   U3080 : NAND4_X1 port map( A1 => n5263, A2 => n5264, A3 => n5265, A4 => 
                           n5262, ZN => n5271);
   U3081 : INV_X1 port map( A => n5266, ZN => n5269);
   U3082 : INV_X1 port map( A => n5267, ZN => n5268);
   U3083 : NAND2_X1 port map( A1 => n5269, A2 => n5268, ZN => n5270);
   U3084 : AND2_X1 port map( A1 => n5271, A2 => n5270, ZN => n7920);
   U3085 : NOR2_X1 port map( A1 => n383, A2 => n365, ZN => n5272);
   U3088 : NAND2_X1 port map( A1 => n5302, A2 => n5273, ZN => n6342);
   U3089 : MUX2_X1 port map( A => n6800, B => n7508, S => n2638, Z => n5276);
   U3090 : XNOR2_X1 port map( A => n8393, B => n6593, ZN => n5274);
   U3091 : NAND2_X1 port map( A1 => n6595, A2 => n5274, ZN => n5275);
   U3092 : NAND2_X1 port map( A1 => n5276, A2 => n5275, ZN => n5480);
   U3093 : XNOR2_X1 port map( A => n371, B => n6259, ZN => n5277);
   U3094 : OAI22_X1 port map( A1 => mult_x_19_n4, A2 => n5277, B1 => n7949, B2 
                           => n8329, ZN => n5481);
   U3095 : XNOR2_X1 port map( A => n5480, B => n5481, ZN => n5279);
   U3096 : MUX2_X1 port map( A => n8500, B => n7053, S => n386, Z => n5479);
   U3097 : NAND2_X1 port map( A1 => n5479, A2 => n5478, ZN => n5278);
   U3098 : XNOR2_X1 port map( A => n5279, B => n5278, ZN => n5460);
   U3099 : AND2_X1 port map( A1 => n5281, A2 => n5280, ZN => n5283);
   U3100 : OAI22_X1 port map( A1 => n5283, A2 => n5282, B1 => n5281, B2 => 
                           n5280, ZN => n5461);
   U3101 : XNOR2_X1 port map( A => n5460, B => n5461, ZN => n5293);
   U3102 : MUX2_X1 port map( A => n8459, B => n8434, S => n4381, Z => n5286);
   U3103 : XNOR2_X1 port map( A => n8326, B => n8002, ZN => n5284);
   U3104 : NAND2_X1 port map( A1 => n6264, A2 => n5284, ZN => n5285);
   U3105 : NAND2_X1 port map( A1 => n5286, A2 => n5285, ZN => n5486);
   U3106 : MUX2_X1 port map( A => n6715, B => n6887, S => n204, Z => n5289);
   U3107 : XNOR2_X1 port map( A => n8392, B => n6244, ZN => n5287);
   U3108 : NAND2_X1 port map( A1 => n7861, A2 => n5287, ZN => n5288);
   U3109 : NAND2_X1 port map( A1 => n5289, A2 => n5288, ZN => n5680);
   U3110 : XNOR2_X1 port map( A => n5486, B => n5680, ZN => n5292);
   U3111 : MUX2_X1 port map( A => n8577, B => n4490, S => B_SIG_9_port, Z => 
                           n5291);
   U3112 : MUX2_X1 port map( A => n8595, B => n4607, S => n6109, Z => n5290);
   U3113 : NAND2_X1 port map( A1 => n5291, A2 => n5290, ZN => n5681);
   U3114 : XNOR2_X1 port map( A => n5293, B => n5470, ZN => n5332);
   U3115 : INV_X1 port map( A => n5332, ZN => n5330);
   U3116 : NAND2_X1 port map( A1 => n5296, A2 => n5297, ZN => n5294);
   U3117 : NAND2_X1 port map( A1 => n5295, A2 => n5294, ZN => n5301);
   U3118 : INV_X1 port map( A => n5296, ZN => n5299);
   U3119 : INV_X1 port map( A => n5297, ZN => n5298);
   U3120 : NAND2_X1 port map( A1 => n5299, A2 => n5298, ZN => n5300);
   U3121 : NAND2_X1 port map( A1 => n5301, A2 => n5300, ZN => n5465);
   U3122 : NAND2_X1 port map( A1 => n8339, A2 => n5508, ZN => n5867);
   U3124 : NAND2_X1 port map( A1 => n7559, A2 => n5303, ZN => n7659);
   U3125 : NAND2_X1 port map( A1 => n7439, A2 => n8354, ZN => n5305);
   U3126 : AND2_X1 port map( A1 => n7659, A2 => n5305, ZN => n5311);
   U3128 : MUX2_X1 port map( A => n7123, B => n7122, S => n390, Z => n5309);
   U3129 : XNOR2_X1 port map( A => n8403, B => n362, ZN => n5306);
   U3130 : NAND2_X1 port map( A1 => n5307, A2 => n5306, ZN => n5308);
   U3131 : NAND2_X1 port map( A1 => n5309, A2 => n5308, ZN => n5310);
   U3132 : NAND2_X1 port map( A1 => n5311, A2 => n5310, ZN => n5421);
   U3133 : INV_X1 port map( A => n5310, ZN => n5313);
   U3134 : INV_X1 port map( A => n5311, ZN => n5312);
   U3135 : NAND2_X1 port map( A1 => n5313, A2 => n5312, ZN => n5314);
   U3136 : NAND2_X1 port map( A1 => n5421, A2 => n5314, ZN => n5466);
   U3137 : XNOR2_X1 port map( A => n5465, B => n5466, ZN => n5328);
   U3138 : OAI22_X1 port map( A1 => n6606, A2 => n7123, B1 => n7122, B2 => 
                           n8401, ZN => n5318);
   U3139 : INV_X1 port map( A => n5315, ZN => n5317);
   U3140 : INV_X1 port map( A => n5324, ZN => n5316);
   U3141 : OAI21_X1 port map( B1 => n5318, B2 => n5317, A => n5316, ZN => n5319
                           );
   U3142 : AND2_X1 port map( A1 => n5320, A2 => n5319, ZN => n5322);
   U3143 : NAND2_X1 port map( A1 => n5322, A2 => n5321, ZN => n5327);
   U3144 : INV_X1 port map( A => n5323, ZN => n5325);
   U3145 : NAND2_X1 port map( A1 => n5325, A2 => n5324, ZN => n5326);
   U3146 : NAND2_X1 port map( A1 => n5327, A2 => n5326, ZN => n5464);
   U3147 : XNOR2_X1 port map( A => n5328, B => n5464, ZN => n5331);
   U3148 : INV_X1 port map( A => n5331, ZN => n5329);
   U3149 : NAND2_X1 port map( A1 => n5330, A2 => n5329, ZN => n5541);
   U3150 : NAND2_X1 port map( A1 => n5332, A2 => n5331, ZN => n5542);
   U3151 : INV_X1 port map( A => n5333, ZN => n5337);
   U3152 : INV_X1 port map( A => n5334, ZN => n5336);
   U3153 : OAI21_X1 port map( B1 => n5337, B2 => n5336, A => n5335, ZN => n5339
                           );
   U3154 : NAND2_X1 port map( A1 => n5337, A2 => n5336, ZN => n5338);
   U3155 : NAND2_X1 port map( A1 => n5339, A2 => n5338, ZN => n5560);
   U3156 : XNOR2_X1 port map( A => n5559, B => n5560, ZN => n5371);
   U3157 : MUX2_X1 port map( A => n7216, B => n7215, S => n6606, Z => n5341);
   U3158 : MUX2_X1 port map( A => n6460, B => n5226, S => n8324, Z => n5340);
   U3159 : NOR2_X2 port map( A1 => n5341, A2 => n5340, ZN => n5677);
   U3160 : MUX2_X1 port map( A => n8488, B => n5395, S => n372, Z => n5343);
   U3161 : MUX2_X1 port map( A => n5398, B => n5397, S => n360, Z => n5342);
   U3162 : NOR2_X1 port map( A1 => n5343, A2 => n5342, ZN => n5674);
   U3163 : NAND2_X1 port map( A1 => n5677, A2 => n5674, ZN => n5492);
   U3164 : NAND2_X1 port map( A1 => n5492, A2 => n5491, ZN => n5346);
   U3165 : MUX2_X1 port map( A => n4975, B => n8012, S => n8332, Z => n5345);
   U3166 : MUX2_X1 port map( A => n8455, B => n8553, S => n359, Z => n5344);
   U3167 : XNOR2_X1 port map( A => n5346, B => n5676, ZN => n5356);
   U3168 : NAND4_X1 port map( A1 => n5350, A2 => n5349, A3 => n5348, A4 => 
                           n5347, ZN => n5355);
   U3169 : NAND3_X1 port map( A1 => n5353, A2 => n5352, A3 => n5351, ZN => 
                           n5354);
   U3170 : AND2_X1 port map( A1 => n5355, A2 => n5354, ZN => n5357);
   U3171 : NAND2_X1 port map( A1 => n5356, A2 => n5357, ZN => n5495);
   U3172 : INV_X1 port map( A => n5356, ZN => n5359);
   U3173 : INV_X1 port map( A => n5357, ZN => n5358);
   U3174 : NAND2_X1 port map( A1 => n5359, A2 => n5358, ZN => n5498);
   U3175 : NAND2_X1 port map( A1 => n5495, A2 => n5498, ZN => n5365);
   U3176 : INV_X1 port map( A => n5360, ZN => n5361);
   U3177 : NAND2_X1 port map( A1 => n5362, A2 => n5361, ZN => n5364);
   U3178 : NAND2_X1 port map( A1 => n5364, A2 => n5363, ZN => n5497);
   U3179 : XNOR2_X1 port map( A => n5365, B => n5497, ZN => n5561);
   U3180 : INV_X1 port map( A => n5366, ZN => n5368);
   U3181 : OAI21_X1 port map( B1 => n5369, B2 => n5368, A => n5367, ZN => n5557
                           );
   U3182 : XNOR2_X1 port map( A => n5561, B => n5557, ZN => n5370);
   U3183 : XNOR2_X1 port map( A => n5371, B => n5370, ZN => n5382);
   U3184 : INV_X1 port map( A => n5376, ZN => n5372);
   U3185 : NAND2_X1 port map( A1 => n4457, A2 => n5372, ZN => n5373);
   U3186 : NAND2_X1 port map( A1 => n5374, A2 => n5373, ZN => n5379);
   U3187 : INV_X1 port map( A => n4457, ZN => n5377);
   U3188 : NAND2_X1 port map( A1 => n5377, A2 => n5376, ZN => n5378);
   U3189 : NAND2_X1 port map( A1 => n5379, A2 => n5378, ZN => n5381);
   U3190 : NAND2_X1 port map( A1 => n5382, A2 => n5381, ZN => n7919);
   U3191 : NAND4_X1 port map( A1 => n7922, A2 => n5380, A3 => n7920, A4 => 
                           n7919, ZN => n8025);
   U3192 : INV_X1 port map( A => n5381, ZN => n5384);
   U3193 : INV_X1 port map( A => n5382, ZN => n5383);
   U3194 : NAND2_X1 port map( A1 => n5384, A2 => n5383, ZN => n8026);
   U3195 : AND2_X1 port map( A1 => n8400, A2 => n8339, ZN => n5385);
   U3197 : AND2_X1 port map( A1 => n370, A2 => n393, ZN => n5386);
   U3198 : BUF_X2 port map( A => n8581, Z => n7695);
   U3199 : MUX2_X1 port map( A => n8559, B => n7695, S => n2638, Z => n5389);
   U3200 : BUF_X2 port map( A => n5407, Z => n6374);
   U3201 : XNOR2_X1 port map( A => n8393, B => n8503, ZN => n5387);
   U3202 : NAND2_X1 port map( A1 => n6374, A2 => n5387, ZN => n5388);
   U3203 : NAND2_X1 port map( A1 => n5389, A2 => n5388, ZN => n5394);
   U3204 : MUX2_X1 port map( A => n7324, B => n7323, S => n8352, Z => n5392);
   U3205 : XNOR2_X1 port map( A => n8369, B => n362, ZN => n5390);
   U3206 : NAND2_X1 port map( A1 => n5041, A2 => n5390, ZN => n5391);
   U3207 : NAND2_X1 port map( A1 => n5392, A2 => n5391, ZN => n5393);
   U3208 : NAND2_X1 port map( A1 => n5394, A2 => n5393, ZN => n5596);
   U3209 : NAND2_X1 port map( A1 => n5598, A2 => n5596, ZN => n5401);
   U3210 : MUX2_X1 port map( A => n8488, B => n5395, S => n371, Z => n5400);
   U3211 : MUX2_X1 port map( A => n5398, B => n5397, S => n363, Z => n5399);
   U3212 : NOR2_X1 port map( A1 => n5400, A2 => n5399, ZN => n5597);
   U3213 : XNOR2_X1 port map( A => n5401, B => n5597, ZN => n5591);
   U3214 : MUX2_X1 port map( A => n7946, B => n7947, S => n205, Z => n5403);
   U3215 : NAND2_X1 port map( A1 => n5781, A2 => n8423, ZN => n5402);
   U3216 : NAND2_X1 port map( A1 => n5403, A2 => n5402, ZN => n5601);
   U3217 : XNOR2_X1 port map( A => n8328, B => n6593, ZN => n5404);
   U3218 : NAND2_X1 port map( A1 => n6595, A2 => n5404, ZN => n5602);
   U3219 : BUF_X2 port map( A => n6800, Z => n7227);
   U3220 : OR2_X1 port map( A1 => n7227, A2 => n381, ZN => n5405);
   U3221 : OAI211_X1 port map( C1 => n7439, C2 => n8396, A => n5602, B => n5405
                           , ZN => n5406);
   U3222 : XNOR2_X1 port map( A => n5601, B => n5406, ZN => n5408);
   U3223 : NOR2_X1 port map( A1 => n8503, A2 => n4430, ZN => n5861);
   U3224 : INV_X1 port map( A => n8582, ZN => n7751);
   U3225 : AOI21_X1 port map( B1 => n7087, B2 => n2638, A => n7751, ZN => n5605
                           );
   U3226 : XNOR2_X1 port map( A => n5408, B => n5605, ZN => n5592);
   U3227 : XNOR2_X1 port map( A => n5591, B => n5592, ZN => n5420);
   U3228 : NAND2_X1 port map( A1 => n5878, A2 => n360, ZN => n5411);
   U3229 : NAND2_X1 port map( A1 => n6102, A2 => n8337, ZN => n5410);
   U3230 : INV_X1 port map( A => n6251, ZN => n6104);
   U3231 : XNOR2_X1 port map( A => n5879, B => n8330, ZN => n5409);
   U3232 : AOI22_X1 port map( A1 => n5411, A2 => n5410, B1 => n6104, B2 => 
                           n5409, ZN => n5652);
   U3233 : XNOR2_X1 port map( A => n5883, B => n8392, ZN => n5412);
   U3234 : NAND2_X1 port map( A1 => n4491, A2 => n5412, ZN => n5414);
   U3235 : NAND3_X1 port map( A1 => n5414, A2 => n204, A3 => n8595, ZN => n5653
                           );
   U3236 : AND2_X1 port map( A1 => n4607, A2 => n8351, ZN => n5413);
   U3237 : NAND2_X1 port map( A1 => n5414, A2 => n5413, ZN => n5654);
   U3238 : NAND2_X1 port map( A1 => n5653, A2 => n5654, ZN => n5415);
   U3239 : NAND2_X1 port map( A1 => n5415, A2 => n5652, ZN => n5658);
   U3240 : OAI21_X1 port map( B1 => n5652, B2 => n5415, A => n5658, ZN => n5419
                           );
   U3241 : INV_X1 port map( A => n4461, ZN => n6362);
   U3242 : INV_X1 port map( A => n7054, ZN => n6361);
   U3243 : MUX2_X1 port map( A => n6362, B => n6361, S => n8350, Z => n5418);
   U3244 : INV_X1 port map( A => n6702, ZN => n6365);
   U3245 : XNOR2_X1 port map( A => n6606, B => n4401, ZN => n5416);
   U3246 : NOR2_X1 port map( A1 => n6365, A2 => n5416, ZN => n5417);
   U3247 : NOR2_X1 port map( A1 => n5418, A2 => n5417, ZN => n5657);
   U3248 : XNOR2_X1 port map( A => n5419, B => n5657, ZN => n5593);
   U3249 : XNOR2_X1 port map( A => n5420, B => n5593, ZN => n5453);
   U3250 : INV_X1 port map( A => n5421, ZN => n5426);
   U3251 : MUX2_X1 port map( A => n8547, B => n8546, S => n360, Z => n5423);
   U3252 : MUX2_X1 port map( A => n5878, B => n6102, S => n8332, Z => n5422);
   U3253 : NAND2_X1 port map( A1 => n5423, A2 => n5422, ZN => n5457);
   U3254 : MUX2_X1 port map( A => n4487, B => n7325, S => n390, Z => n5425);
   U3255 : MUX2_X1 port map( A => n7324, B => n8465, S => n8401, Z => n5424);
   U3256 : NAND2_X1 port map( A1 => n5425, A2 => n5424, ZN => n5456);
   U3257 : OAI21_X1 port map( B1 => n5426, B2 => n5457, A => n5456, ZN => n5428
                           );
   U3258 : NAND2_X1 port map( A1 => n5426, A2 => n5457, ZN => n5427);
   U3259 : NAND2_X1 port map( A1 => n5428, A2 => n5427, ZN => n5583);
   U3260 : MUX2_X1 port map( A => n6362, B => n6361, S => n8328, Z => n5431);
   U3261 : XNOR2_X1 port map( A => n4401, B => n8324, ZN => n5429);
   U3262 : NOR2_X1 port map( A1 => n6365, A2 => n5429, ZN => n5430);
   U3263 : NOR2_X1 port map( A1 => n5431, A2 => n5430, ZN => n5439);
   U3264 : INV_X1 port map( A => n7947, ZN => n5433);
   U3265 : INV_X1 port map( A => n7946, ZN => n5432);
   U3267 : NOR2_X1 port map( A1 => n7949, A2 => n8325, ZN => n5434);
   U3269 : INV_X1 port map( A => n5440, ZN => n5436);
   U3270 : NAND2_X1 port map( A1 => n4460, A2 => n5436, ZN => n5499);
   U3271 : INV_X1 port map( A => n5499, ZN => n5441);
   U3272 : MUX2_X1 port map( A => n8445, B => n6740, S => n359, Z => n5438);
   U3273 : MUX2_X1 port map( A => n8459, B => n8434, S => n8326, Z => n5437);
   U3274 : NAND2_X1 port map( A1 => n5438, A2 => n5437, ZN => n5501);
   U3275 : NAND2_X1 port map( A1 => n5439, A2 => n5440, ZN => n5500);
   U3276 : MUX2_X1 port map( A => n5898, B => n6249, S => n363, Z => n5443);
   U3277 : MUX2_X1 port map( A => n8454, B => n8515, S => n372, Z => n5442);
   U3278 : NAND2_X1 port map( A1 => n5443, A2 => n5442, ZN => n5513);
   U3279 : INV_X1 port map( A => n5513, ZN => n5451);
   U3280 : MUX2_X1 port map( A => n4489, B => n8577, S => n204, Z => n5445);
   U3281 : MUX2_X1 port map( A => n4607, B => n8596, S => n8327, Z => n5444);
   U3282 : NAND2_X1 port map( A1 => n5445, A2 => n5444, ZN => n5514);
   U3283 : XNOR2_X1 port map( A => n4381, B => n6244, ZN => n5446);
   U3284 : NAND2_X1 port map( A1 => n7861, A2 => n5446, ZN => n5447);
   U3285 : NAND2_X1 port map( A1 => n5514, A2 => n5512, ZN => n5450);
   U3286 : INV_X1 port map( A => n5514, ZN => n5449);
   U3287 : INV_X1 port map( A => n5512, ZN => n5448);
   U3289 : NAND2_X1 port map( A1 => n5453, A2 => n5452, ZN => n5581);
   U3290 : NAND2_X1 port map( A1 => n5581, A2 => n5580, ZN => n5476);
   U3291 : INV_X1 port map( A => n5461, ZN => n5454);
   U3292 : NAND2_X1 port map( A1 => n5460, A2 => n5454, ZN => n5474);
   U3293 : INV_X1 port map( A => n5470, ZN => n5455);
   U3294 : NAND2_X1 port map( A1 => n5474, A2 => n5455, ZN => n5463);
   U3295 : XNOR2_X1 port map( A => n5421, B => n5456, ZN => n5459);
   U3296 : INV_X1 port map( A => n5457, ZN => n5458);
   U3297 : XNOR2_X1 port map( A => n5459, B => n5458, ZN => n5472);
   U3299 : NAND2_X1 port map( A1 => n8495, A2 => n5461, ZN => n5471);
   U3300 : AND3_X1 port map( A1 => n5463, A2 => n5472, A3 => n5471, ZN => n5545
                           );
   U3301 : INV_X1 port map( A => n5464, ZN => n5469);
   U3302 : INV_X1 port map( A => n5465, ZN => n5468);
   U3303 : INV_X1 port map( A => n5466, ZN => n5467);
   U3304 : FA_X1 port map( A => n5469, B => n5468, CI => n5467, CO => n5547, S 
                           => n_1134);
   U3305 : NAND2_X1 port map( A1 => n5471, A2 => n5470, ZN => n5475);
   U3306 : INV_X1 port map( A => n5472, ZN => n5473);
   U3307 : NAND3_X1 port map( A1 => n5475, A2 => n5474, A3 => n5473, ZN => 
                           n5544);
   U3308 : OAI21_X1 port map( B1 => n5545, B2 => n5547, A => n5544, ZN => n5579
                           );
   U3309 : XNOR2_X1 port map( A => n5476, B => n5579, ZN => n5830);
   U3310 : AND2_X1 port map( A1 => n5486, A2 => n5680, ZN => n5488);
   U3311 : NAND2_X1 port map( A1 => n8533, A2 => n5481, ZN => n5477);
   U3312 : NAND3_X1 port map( A1 => n5479, A2 => n5478, A3 => n5477, ZN => 
                           n5485);
   U3313 : INV_X1 port map( A => n5480, ZN => n5483);
   U3314 : INV_X1 port map( A => n5481, ZN => n5482);
   U3315 : NAND2_X1 port map( A1 => n5483, A2 => n5482, ZN => n5484);
   U3316 : INV_X1 port map( A => n5486, ZN => n5682);
   U3317 : INV_X1 port map( A => n5680, ZN => n5684);
   U3318 : NAND2_X1 port map( A1 => n5682, A2 => n5684, ZN => n5487);
   U3319 : OAI211_X1 port map( C1 => n5488, C2 => n5681, A => n5678, B => n5487
                           , ZN => n5530);
   U3320 : INV_X1 port map( A => n5681, ZN => n5685);
   U3321 : INV_X1 port map( A => n5487, ZN => n5490);
   U3322 : INV_X1 port map( A => n5678, ZN => n5670);
   U3323 : INV_X1 port map( A => n5488, ZN => n5489);
   U3324 : OAI211_X1 port map( C1 => n5685, C2 => n5490, A => n5670, B => n5489
                           , ZN => n5531);
   U3325 : NAND2_X1 port map( A1 => n5530, A2 => n5531, ZN => n5494);
   U3326 : NAND2_X1 port map( A1 => n5491, A2 => n5676, ZN => n5493);
   U3327 : XNOR2_X1 port map( A => n5494, B => n5669, ZN => n5551);
   U3328 : INV_X1 port map( A => n5495, ZN => n5496);
   U3329 : NAND2_X1 port map( A1 => n5500, A2 => n5499, ZN => n5502);
   U3330 : XNOR2_X1 port map( A => n5502, B => n5501, ZN => n5534);
   U3331 : INV_X1 port map( A => n7120, ZN => n7232);
   U3332 : MUX2_X1 port map( A => n7232, B => n7012, S => n6109, Z => n5505);
   U3333 : INV_X1 port map( A => n8593, ZN => n7231);
   U3334 : MUX2_X1 port map( A => n7231, B => n7010, S => n362, Z => n5504);
   U3335 : NOR2_X1 port map( A1 => n5505, A2 => n5504, ZN => n5507);
   U3336 : NAND2_X1 port map( A1 => n6374, A2 => n8354, ZN => n5506);
   U3337 : NAND2_X1 port map( A1 => n5507, A2 => n5506, ZN => n5524);
   U3338 : NAND2_X1 port map( A1 => n5524, A2 => n5526, ZN => n5511);
   U3339 : MUX2_X1 port map( A => n8476, B => n7559, S => n381, Z => n5510);
   U3340 : MUX2_X1 port map( A => n7227, B => n7439, S => n395, Z => n5509);
   U3341 : NAND2_X1 port map( A1 => n5510, A2 => n5509, ZN => n5525);
   U3342 : XNOR2_X1 port map( A => n5511, B => n5525, ZN => n5536);
   U3343 : XNOR2_X1 port map( A => n5536, B => n5534, ZN => n5549);
   U3344 : XNOR2_X1 port map( A => n5513, B => n5512, ZN => n5515);
   U3345 : XNOR2_X1 port map( A => n5549, B => n5553, ZN => n5516);
   U3346 : MUX2_X1 port map( A => n7120, B => n7121, S => B_SIG_9_port, Z => 
                           n5518);
   U3347 : MUX2_X1 port map( A => n6812, B => n7123, S => n7945, Z => n5517);
   U3348 : NAND2_X1 port map( A1 => n5518, A2 => n5517, ZN => n5772);
   U3349 : MUX2_X1 port map( A => n6715, B => n6887, S => n373, Z => n5521);
   U3350 : XNOR2_X1 port map( A => n8326, B => n6244, ZN => n5519);
   U3351 : NAND2_X1 port map( A1 => n7861, A2 => n5519, ZN => n5520);
   U3352 : NAND2_X1 port map( A1 => n5521, A2 => n5520, ZN => n5641);
   U3353 : XNOR2_X1 port map( A => n5772, B => n5641, ZN => n5523);
   U3354 : MUX2_X1 port map( A => n8445, B => n6740, S => n377, Z => n5639);
   U3355 : MUX2_X1 port map( A => n8459, B => n8434, S => n8394, Z => n5636);
   U3356 : XNOR2_X1 port map( A => n5523, B => n5522, ZN => n5529);
   U3357 : INV_X1 port map( A => n5524, ZN => n5528);
   U3358 : INV_X1 port map( A => n5525, ZN => n5527);
   U3359 : OAI21_X1 port map( B1 => n5528, B2 => n5527, A => n5526, ZN => n5644
                           );
   U3360 : XNOR2_X1 port map( A => n5529, B => n5644, ZN => n5690);
   U3361 : INV_X1 port map( A => n5530, ZN => n5532);
   U3362 : OAI21_X1 port map( B1 => n5532, B2 => n5669, A => n8539, ZN => n5533
                           );
   U3363 : XNOR2_X1 port map( A => n5690, B => n5533, ZN => n5540);
   U3364 : NAND2_X1 port map( A1 => n5536, A2 => n5553, ZN => n5699);
   U3365 : INV_X1 port map( A => n5534, ZN => n5535);
   U3366 : NAND2_X1 port map( A1 => n5699, A2 => n5535, ZN => n5689);
   U3367 : INV_X1 port map( A => n5536, ZN => n5538);
   U3368 : INV_X1 port map( A => n5553, ZN => n5537);
   U3369 : NAND2_X1 port map( A1 => n5538, A2 => n5537, ZN => n5693);
   U3370 : NAND2_X1 port map( A1 => n5689, A2 => n5693, ZN => n5539);
   U3371 : NAND2_X1 port map( A1 => n5541, A2 => n5557, ZN => n5543);
   U3372 : INV_X1 port map( A => n5544, ZN => n5546);
   U3373 : XNOR2_X1 port map( A => n5548, B => n5547, ZN => n5566);
   U3374 : XNOR2_X1 port map( A => n8431, B => n5549, ZN => n5555);
   U3377 : XNOR2_X1 port map( A => n5554, B => n5555, ZN => n5565);
   U3378 : FA_X1 port map( A => n5568, B => n5566, CI => n5565, CO => n5575, S 
                           => n_1135);
   U3380 : XNOR2_X1 port map( A => n8496, B => n5568, ZN => n5569);
   U3381 : XNOR2_X1 port map( A => n4504, B => n5569, ZN => n5572);
   U3383 : INV_X1 port map( A => n5571, ZN => n5574);
   U3384 : NAND2_X1 port map( A1 => n5572, A2 => n5573, ZN => n5577);
   U3385 : NAND2_X1 port map( A1 => n5577, A2 => n5574, ZN => n5576);
   U3386 : NAND2_X1 port map( A1 => n5576, A2 => n5575, ZN => n7933);
   U3387 : INV_X1 port map( A => n5577, ZN => n5578);
   U3388 : NAND2_X1 port map( A1 => n5571, A2 => n5578, ZN => n7934);
   U3389 : NAND2_X1 port map( A1 => n5580, A2 => n5579, ZN => n5582);
   U3390 : NAND2_X1 port map( A1 => n5582, A2 => n5581, ZN => n5824);
   U3391 : NAND2_X1 port map( A1 => n5586, A2 => n5583, ZN => n5585);
   U3392 : NAND2_X1 port map( A1 => n5585, A2 => n5584, ZN => n5590);
   U3393 : INV_X1 port map( A => n5583, ZN => n5588);
   U3394 : INV_X1 port map( A => n5586, ZN => n5587);
   U3395 : NAND2_X1 port map( A1 => n5588, A2 => n5587, ZN => n5589);
   U3396 : NAND2_X1 port map( A1 => n5590, A2 => n5589, ZN => n5814);
   U3397 : OAI21_X1 port map( B1 => n5593, B2 => n8583, A => n5592, ZN => n5595
                           );
   U3398 : NAND2_X1 port map( A1 => n5593, A2 => n8583, ZN => n5594);
   U3399 : NAND2_X1 port map( A1 => n5595, A2 => n5594, ZN => n5815);
   U3400 : XNOR2_X1 port map( A => n5814, B => n5815, ZN => n5609);
   U3401 : INV_X1 port map( A => n5596, ZN => n5600);
   U3402 : INV_X1 port map( A => n5597, ZN => n5599);
   U3403 : OAI21_X1 port map( B1 => n5600, B2 => n5599, A => n5598, ZN => n5811
                           );
   U3404 : INV_X1 port map( A => n5601, ZN => n5604);
   U3405 : MUX2_X1 port map( A => n8568, B => n7439, S => n381, Z => n5603);
   U3406 : OAI211_X1 port map( C1 => n5605, C2 => n5604, A => n5603, B => n5602
                           , ZN => n5607);
   U3407 : NAND2_X1 port map( A1 => n5605, A2 => n5604, ZN => n5606);
   U3408 : NAND2_X1 port map( A1 => n5607, A2 => n5606, ZN => n5774);
   U3409 : XNOR2_X1 port map( A => n5811, B => n5774, ZN => n5608);
   U3410 : NAND2_X1 port map( A1 => n5771, A2 => n5772, ZN => n5810);
   U3411 : XNOR2_X1 port map( A => n5608, B => n5810, ZN => n5816);
   U3412 : XNOR2_X1 port map( A => n5609, B => n5816, ZN => n5823);
   U3413 : MUX2_X1 port map( A => n5898, B => n6249, S => n8423, Z => n5611);
   U3414 : MUX2_X1 port map( A => n6126, B => n6248, S => n371, Z => n5610);
   U3415 : NAND2_X1 port map( A1 => n5611, A2 => n5610, ZN => n5789);
   U3416 : MUX2_X1 port map( A => n4490, B => n7051, S => n373, Z => n5613);
   U3417 : MUX2_X1 port map( A => n4607, B => n8596, S => n379, Z => n5612);
   U3418 : NAND2_X1 port map( A1 => n5613, A2 => n5612, ZN => n5785);
   U3419 : XNOR2_X1 port map( A => n5789, B => n5785, ZN => n5616);
   U3420 : MUX2_X1 port map( A => n8501, B => n7053, S => n390, Z => n5615);
   U3421 : MUX2_X1 port map( A => n4462, B => n7198, S => n8401, Z => n5614);
   U3422 : NAND2_X1 port map( A1 => n5615, A2 => n5614, ZN => n5788);
   U3423 : XNOR2_X1 port map( A => n5616, B => n5788, ZN => n5631);
   U3424 : INV_X1 port map( A => n6819, ZN => n5873);
   U3425 : MUX2_X1 port map( A => n5873, B => n5872, S => n356, Z => n5619);
   U3426 : INV_X1 port map( A => n7861, ZN => n5875);
   U3427 : XNOR2_X1 port map( A => n359, B => n6244, ZN => n5617);
   U3428 : NOR2_X1 port map( A1 => n5875, A2 => n5617, ZN => n5618);
   U3429 : MUX2_X1 port map( A => n7324, B => n7323, S => n8333, Z => n5623);
   U3431 : XNOR2_X1 port map( A => n6229, B => n7945, ZN => n5621);
   U3432 : NAND2_X1 port map( A1 => n5621, A2 => n5041, ZN => n5622);
   U3433 : INV_X1 port map( A => n5626, ZN => n5624);
   U3434 : NAND2_X1 port map( A1 => n5625, A2 => n5624, ZN => n5716);
   U3435 : NAND2_X1 port map( A1 => n5627, A2 => n5626, ZN => n5714);
   U3436 : NAND2_X1 port map( A1 => n5716, A2 => n5714, ZN => n5630);
   U3437 : MUX2_X1 port map( A => n5845, B => n5844, S => n363, Z => n5629);
   U3438 : MUX2_X1 port map( A => n6103, B => n6102, S => n8330, Z => n5628);
   U3439 : NAND2_X1 port map( A1 => n5629, A2 => n5628, ZN => n5713);
   U3440 : XNOR2_X1 port map( A => n5630, B => n5713, ZN => n5632);
   U3441 : NAND2_X1 port map( A1 => n5631, A2 => n5632, ZN => n5972);
   U3442 : INV_X1 port map( A => n5631, ZN => n5634);
   U3443 : INV_X1 port map( A => n5632, ZN => n5633);
   U3444 : NAND2_X1 port map( A1 => n5634, A2 => n5633, ZN => n5732);
   U3445 : NAND2_X1 port map( A1 => n5972, A2 => n5732, ZN => n5645);
   U3446 : INV_X1 port map( A => n5772, ZN => n5640);
   U3447 : INV_X1 port map( A => n5636, ZN => n5635);
   U3448 : AOI21_X1 port map( B1 => n5640, B2 => n5635, A => n5641, ZN => n5638
                           );
   U3449 : NAND3_X1 port map( A1 => n5772, A2 => n5639, A3 => n5636, ZN => 
                           n5637);
   U3450 : OAI211_X1 port map( C1 => n5639, C2 => n5772, A => n5638, B => n5637
                           , ZN => n5643);
   U3451 : XNOR2_X1 port map( A => n5771, B => n5640, ZN => n5642);
   U3453 : XNOR2_X1 port map( A => n5645, B => n5968, ZN => n5706);
   U3454 : XNOR2_X1 port map( A => n8350, B => n6593, ZN => n5646);
   U3455 : NAND2_X1 port map( A1 => n6595, A2 => n5646, ZN => n5647);
   U3456 : XNOR2_X1 port map( A => n6113, B => n200, ZN => n5744);
   U3457 : INV_X1 port map( A => n5749, ZN => n5648);
   U3458 : NOR2_X1 port map( A1 => n5648, A2 => n2638, ZN => n5722);
   U3459 : XNOR2_X1 port map( A => n8556, B => n5722, ZN => n5651);
   U3460 : MUX2_X1 port map( A => n7123, B => n7122, S => n8327, Z => n5649);
   U3461 : NAND2_X1 port map( A1 => n5650, A2 => n5649, ZN => n5718);
   U3462 : XNOR2_X1 port map( A => n5651, B => n5718, ZN => n5707);
   U3463 : INV_X1 port map( A => n5652, ZN => n5655);
   U3464 : NAND3_X1 port map( A1 => n5655, A2 => n5654, A3 => n5653, ZN => 
                           n5656);
   U3465 : NAND2_X1 port map( A1 => n5657, A2 => n5656, ZN => n5659);
   U3466 : NAND2_X1 port map( A1 => n5659, A2 => n5658, ZN => n5711);
   U3467 : XNOR2_X1 port map( A => n5707, B => n5711, ZN => n5668);
   U3468 : MUX2_X1 port map( A => n7696, B => n7695, S => n395, Z => n5662);
   U3469 : XNOR2_X1 port map( A => n8396, B => n8503, ZN => n5660);
   U3470 : NAND2_X1 port map( A1 => n6374, A2 => n5660, ZN => n5661);
   U3471 : NAND2_X1 port map( A1 => n5662, A2 => n5661, ZN => n5728);
   U3472 : MUX2_X1 port map( A => n7946, B => n7947, S => n357, Z => n5664);
   U3473 : NAND2_X1 port map( A1 => n5781, A2 => n205, ZN => n5663);
   U3474 : NAND2_X1 port map( A1 => n5664, A2 => n5663, ZN => n5727);
   U3475 : XNOR2_X1 port map( A => n5728, B => n5727, ZN => n5667);
   U3476 : MUX2_X1 port map( A => n8445, B => n6740, S => n360, Z => n5666);
   U3477 : MUX2_X1 port map( A => n8459, B => n8434, S => n8332, Z => n5665);
   U3478 : NAND2_X1 port map( A1 => n5666, A2 => n5665, ZN => n5730);
   U3479 : XNOR2_X1 port map( A => n5667, B => n5730, ZN => n5708);
   U3480 : XNOR2_X1 port map( A => n5668, B => n5708, ZN => n5705);
   U3481 : XNOR2_X1 port map( A => n8544, B => n5705, ZN => n5703);
   U3482 : INV_X1 port map( A => n5669, ZN => n5671);
   U3483 : NAND2_X1 port map( A1 => n5671, A2 => n5670, ZN => n5696);
   U3484 : INV_X1 port map( A => n5676, ZN => n5673);
   U3485 : INV_X1 port map( A => n5677, ZN => n5672);
   U3486 : NAND2_X1 port map( A1 => n5673, A2 => n5672, ZN => n5675);
   U3487 : AOI22_X1 port map( A1 => n5677, A2 => n5676, B1 => n5675, B2 => 
                           n5674, ZN => n5679);
   U3488 : NAND2_X1 port map( A1 => n5679, A2 => n5678, ZN => n5697);
   U3489 : NAND2_X1 port map( A1 => n5681, A2 => n5680, ZN => n5683);
   U3490 : NAND2_X1 port map( A1 => n5683, A2 => n5682, ZN => n5687);
   U3491 : NAND2_X1 port map( A1 => n5685, A2 => n5684, ZN => n5686);
   U3492 : NAND2_X1 port map( A1 => n5687, A2 => n5686, ZN => n5694);
   U3493 : NAND2_X1 port map( A1 => n5697, A2 => n5694, ZN => n5688);
   U3494 : NAND4_X1 port map( A1 => n5689, A2 => n5693, A3 => n5696, A4 => 
                           n5688, ZN => n5692);
   U3495 : INV_X1 port map( A => n5690, ZN => n5691);
   U3496 : NAND2_X1 port map( A1 => n5692, A2 => n5691, ZN => n5702);
   U3497 : NAND2_X1 port map( A1 => n5693, A2 => n5534, ZN => n5700);
   U3498 : INV_X1 port map( A => n5694, ZN => n5695);
   U3499 : NAND2_X1 port map( A1 => n5696, A2 => n5695, ZN => n5698);
   U3500 : NAND4_X1 port map( A1 => n5700, A2 => n5699, A3 => n5698, A4 => 
                           n5697, ZN => n5701);
   U3501 : NAND2_X1 port map( A1 => n5702, A2 => n5701, ZN => n5704);
   U3502 : XNOR2_X1 port map( A => n5703, B => n5704, ZN => n5822);
   U3503 : FA_X1 port map( A => n5824, B => n5823, CI => n5822, CO => n6064, S 
                           => n_1136);
   U3504 : NAND2_X1 port map( A1 => n8544, A2 => n5705, ZN => n6068);
   U3505 : NAND2_X1 port map( A1 => n6071, A2 => n6068, ZN => n5736);
   U3506 : NAND2_X1 port map( A1 => n5707, A2 => n5708, ZN => n5712);
   U3507 : INV_X1 port map( A => n5707, ZN => n5710);
   U3508 : INV_X1 port map( A => n5708, ZN => n5709);
   U3509 : AOI22_X1 port map( A1 => n5712, A2 => n5711, B1 => n5710, B2 => 
                           n5709, ZN => n5970);
   U3510 : INV_X1 port map( A => n5713, ZN => n5715);
   U3511 : NAND2_X1 port map( A1 => n5715, A2 => n5714, ZN => n5717);
   U3512 : NAND2_X1 port map( A1 => n5717, A2 => n5716, ZN => n5957);
   U3513 : INV_X1 port map( A => n5718, ZN => n5720);
   U3514 : NAND2_X1 port map( A1 => n5721, A2 => n5722, ZN => n5719);
   U3515 : NAND2_X1 port map( A1 => n5720, A2 => n5719, ZN => n5726);
   U3516 : INV_X1 port map( A => n8556, ZN => n5724);
   U3517 : INV_X1 port map( A => n5722, ZN => n5723);
   U3518 : NAND2_X1 port map( A1 => n5724, A2 => n5723, ZN => n5725);
   U3519 : NAND2_X1 port map( A1 => n5726, A2 => n5725, ZN => n5958);
   U3520 : XNOR2_X1 port map( A => n5957, B => n5958, ZN => n5731);
   U3521 : AND2_X1 port map( A1 => n5728, A2 => n5727, ZN => n5729);
   U3522 : OAI22_X1 port map( A1 => n5730, A2 => n5729, B1 => n5728, B2 => 
                           n5727, ZN => n5959);
   U3523 : XNOR2_X1 port map( A => n5731, B => n5959, ZN => n5971);
   U3524 : XNOR2_X1 port map( A => n5970, B => n5971, ZN => n5735);
   U3525 : INV_X1 port map( A => n5732, ZN => n5733);
   U3526 : AOI21_X1 port map( B1 => n5968, B2 => n5972, A => n5733, ZN => n5734
                           );
   U3527 : XNOR2_X1 port map( A => n5736, B => n6073, ZN => n5821);
   U3528 : MUX2_X1 port map( A => n5898, B => n6249, S => n205, Z => n5738);
   U3529 : MUX2_X1 port map( A => n6126, B => n8515, S => n8423, Z => n5737);
   U3530 : NAND2_X1 port map( A1 => n5738, A2 => n5737, ZN => n6013);
   U3531 : MUX2_X1 port map( A => n4462, B => n7198, S => n8352, Z => n5741);
   U3532 : XNOR2_X1 port map( A => n8353, B => n362, ZN => n5739);
   U3533 : NAND2_X1 port map( A1 => n6702, A2 => n5739, ZN => n5740);
   U3534 : NAND2_X1 port map( A1 => n5741, A2 => n5740, ZN => n6012);
   U3535 : XNOR2_X1 port map( A => n6013, B => n6012, ZN => n5767);
   U3536 : MUX2_X1 port map( A => n4489, B => n8577, S => n356, Z => n5743);
   U3537 : MUX2_X1 port map( A => n4607, B => n8596, S => n373, Z => n5742);
   U3538 : AND2_X1 port map( A1 => n5743, A2 => n5742, ZN => n6011);
   U3539 : XNOR2_X1 port map( A => n6011, B => n5767, ZN => n5766);
   U3540 : AND2_X2 port map( A1 => n5744, A2 => n8504, ZN => n7690);
   U3541 : NAND2_X1 port map( A1 => n200, A2 => n387, ZN => n5747);
   U3542 : INV_X1 port map( A => n5747, ZN => n5745);
   U3543 : NAND2_X2 port map( A1 => n5745, A2 => A_SIG_23_port, ZN => n7692);
   U3544 : AOI21_X1 port map( B1 => n7690, B2 => n2638, A => n5746, ZN => n5753
                           );
   U3545 : OAI21_X1 port map( B1 => n5747, B2 => n8354, A => n8504, ZN => n5752
                           );
   U3546 : OAI21_X1 port map( B1 => n5748, B2 => n2638, A => n8398, ZN => n5751
                           );
   U3547 : XNOR2_X1 port map( A => A_SIG_23_port, B => n395, ZN => n5750);
   U3548 : AOI22_X1 port map( A1 => n5752, A2 => n5751, B1 => n5750, B2 => 
                           n5749, ZN => n5754);
   U3549 : NAND2_X1 port map( A1 => n5753, A2 => n5754, ZN => n5924);
   U3550 : INV_X1 port map( A => n5753, ZN => n5756);
   U3551 : INV_X1 port map( A => n5754, ZN => n5755);
   U3552 : NAND2_X1 port map( A1 => n5756, A2 => n5755, ZN => n5926);
   U3553 : NAND2_X1 port map( A1 => n5924, A2 => n5926, ZN => n5765);
   U3554 : MUX2_X1 port map( A => n6800, B => n7439, S => n8324, Z => n5759);
   U3555 : XNOR2_X1 port map( A => n8401, B => n6593, ZN => n5757);
   U3556 : NAND2_X1 port map( A1 => n6595, A2 => n5757, ZN => n5758);
   U3557 : NAND2_X1 port map( A1 => n5759, A2 => n5758, ZN => n5935);
   U3558 : INV_X1 port map( A => n6264, ZN => n8007);
   U3559 : XNOR2_X1 port map( A => n372, B => n8002, ZN => n5764);
   U3560 : INV_X1 port map( A => n6738, ZN => n6743);
   U3561 : OAI21_X1 port map( B1 => n6743, B2 => n8337, A => n5879, ZN => n5762
                           );
   U3562 : OAI21_X1 port map( B1 => n5760, B2 => n360, A => n8397, ZN => n5761)
                           ;
   U3563 : NAND2_X1 port map( A1 => n5762, A2 => n5761, ZN => n5763);
   U3564 : OAI21_X1 port map( B1 => n8007, B2 => n5764, A => n5763, ZN => n5934
                           );
   U3565 : XNOR2_X1 port map( A => n5935, B => n5934, ZN => n5923);
   U3566 : XNOR2_X1 port map( A => n5765, B => n5923, ZN => n5768);
   U3567 : NAND2_X1 port map( A1 => n5766, A2 => n5768, ZN => n6047);
   U3568 : XOR2_X1 port map( A => n5767, B => n6011, Z => n5770);
   U3569 : INV_X1 port map( A => n5768, ZN => n5769);
   U3570 : NAND2_X1 port map( A1 => n5770, A2 => n5769, ZN => n6046);
   U3571 : NAND2_X1 port map( A1 => n6047, A2 => n6046, ZN => n5776);
   U3572 : NAND3_X1 port map( A1 => n4415, A2 => n5772, A3 => n5771, ZN => 
                           n5773);
   U3573 : NAND2_X1 port map( A1 => n5773, A2 => n5811, ZN => n5775);
   U3574 : NAND2_X1 port map( A1 => n5810, A2 => n5774, ZN => n5809);
   U3575 : NAND2_X1 port map( A1 => n5775, A2 => n5809, ZN => n6045);
   U3576 : XNOR2_X1 port map( A => n5776, B => n6045, ZN => n5808);
   U3577 : MUX2_X1 port map( A => n8559, B => n8582, S => n381, Z => n5780);
   U3579 : XNOR2_X1 port map( A => n8328, B => n8503, ZN => n5778);
   U3580 : NAND2_X1 port map( A1 => n6374, A2 => n5778, ZN => n5779);
   U3581 : NAND2_X1 port map( A1 => n5780, A2 => n5779, ZN => n5947);
   U3583 : MUX2_X1 port map( A => n7946, B => n7947, S => n7769, Z => n5783);
   U3584 : NAND2_X1 port map( A1 => n5781, A2 => n357, ZN => n5782);
   U3585 : NAND2_X1 port map( A1 => n5783, A2 => n5782, ZN => n5941);
   U3586 : XNOR2_X1 port map( A => n5947, B => n5941, ZN => n5784);
   U3587 : MUX2_X1 port map( A => n8593, B => n7122, S => n204, Z => n5940);
   U3588 : NAND2_X1 port map( A1 => n5945, A2 => n5940, ZN => n5948);
   U3589 : XNOR2_X1 port map( A => n5784, B => n5948, ZN => n6041);
   U3590 : NAND2_X1 port map( A1 => n5788, A2 => n5789, ZN => n5787);
   U3591 : INV_X1 port map( A => n5785, ZN => n5786);
   U3592 : NAND2_X1 port map( A1 => n5787, A2 => n5786, ZN => n5792);
   U3593 : INV_X1 port map( A => n5788, ZN => n5790);
   U3594 : NAND2_X1 port map( A1 => n5790, A2 => n4458, ZN => n5791);
   U3595 : NAND2_X1 port map( A1 => n5792, A2 => n5791, ZN => n6038);
   U3596 : XNOR2_X1 port map( A => n6041, B => n6038, ZN => n5806);
   U3597 : MUX2_X1 port map( A => n4975, B => n8012, S => n8325, Z => n5796);
   U3598 : MUX2_X1 port map( A => n8455, B => n8553, S => n363, Z => n5795);
   U3599 : NOR2_X1 port map( A1 => n5796, A2 => n5795, ZN => n5799);
   U3600 : MUX2_X1 port map( A => n7215, B => n7216, S => B_SIG_9_port, Z => 
                           n5798);
   U3601 : MUX2_X1 port map( A => n5226, B => n6460, S => n6109, Z => n5797);
   U3602 : NOR2_X1 port map( A1 => n5798, A2 => n5797, ZN => n5800);
   U3603 : NAND2_X1 port map( A1 => n5799, A2 => n5800, ZN => n6020);
   U3604 : INV_X1 port map( A => n5799, ZN => n5802);
   U3605 : INV_X1 port map( A => n5800, ZN => n5801);
   U3606 : NAND2_X1 port map( A1 => n5802, A2 => n5801, ZN => n6019);
   U3607 : NAND2_X1 port map( A1 => n6020, A2 => n6019, ZN => n5805);
   U3608 : MUX2_X1 port map( A => n6714, B => n6888, S => n377, Z => n5804);
   U3609 : MUX2_X1 port map( A => n6715, B => n6887, S => n359, Z => n5803);
   U3610 : NAND2_X1 port map( A1 => n5804, A2 => n5803, ZN => n6017);
   U3611 : XNOR2_X1 port map( A => n5805, B => n6017, ZN => n6040);
   U3612 : XNOR2_X1 port map( A => n5806, B => n6040, ZN => n5807);
   U3613 : NAND2_X1 port map( A1 => n5808, A2 => n5807, ZN => n6056);
   U3614 : NAND2_X1 port map( A1 => n6056, A2 => n6054, ZN => n5820);
   U3615 : INV_X1 port map( A => n5815, ZN => n5819);
   U3616 : OAI21_X1 port map( B1 => n5774, B2 => n5810, A => n5809, ZN => n5813
                           );
   U3617 : INV_X1 port map( A => n5811, ZN => n5812);
   U3618 : XNOR2_X1 port map( A => n5813, B => n5812, ZN => n5818);
   U3619 : OAI21_X1 port map( B1 => n5816, B2 => n5815, A => n5814, ZN => n5817
                           );
   U3620 : OAI21_X1 port map( B1 => n5819, B2 => n5818, A => n5817, ZN => n6055
                           );
   U3621 : XNOR2_X1 port map( A => n5821, B => n8540, ZN => n6065);
   U3622 : NAND2_X1 port map( A1 => n6065, A2 => n6064, ZN => n8033);
   U3623 : INV_X1 port map( A => n5822, ZN => n5826);
   U3624 : XNOR2_X1 port map( A => n5824, B => n5823, ZN => n5825);
   U3626 : INV_X1 port map( A => n5827, ZN => n5831);
   U3627 : INV_X1 port map( A => n5828, ZN => n5829);
   U3628 : FA_X1 port map( A => n5831, B => n5830, CI => n5829, CO => n5833, S 
                           => n_1137);
   U3629 : NAND2_X1 port map( A1 => n8492, A2 => n5833, ZN => n7935);
   U3630 : NAND4_X1 port map( A1 => n7933, A2 => n7934, A3 => n8033, A4 => 
                           n7935, ZN => n6087);
   U3631 : INV_X1 port map( A => n5833, ZN => n8036);
   U3632 : NAND2_X1 port map( A1 => n8033, A2 => n8031, ZN => n6085);
   U3633 : MUX2_X1 port map( A => n6126, B => n6248, S => n357, Z => n5837);
   U3634 : XNOR2_X1 port map( A => n8356, B => n7506, ZN => n5834);
   U3635 : NAND2_X1 port map( A1 => n5835, A2 => n5834, ZN => n5836);
   U3638 : XNOR2_X1 port map( A => B_SIG_9_port, B => n6363, ZN => n5838);
   U3639 : NAND2_X1 port map( A1 => n6702, A2 => n5838, ZN => n5839);
   U3640 : NAND2_X1 port map( A1 => n5840, A2 => n5839, ZN => n6152);
   U3641 : XNOR2_X1 port map( A => n6152, B => n6153, ZN => n5843);
   U3642 : MUX2_X1 port map( A => n7195, B => n7080, S => n379, Z => n5842);
   U3643 : MUX2_X1 port map( A => n7324, B => n8465, S => n8351, Z => n5841);
   U3644 : NAND2_X1 port map( A1 => n5842, A2 => n5841, ZN => n6149);
   U3645 : XNOR2_X1 port map( A => n5843, B => n6149, ZN => n6136);
   U3646 : MUX2_X1 port map( A => n5845, B => n5844, S => n205, Z => n5853);
   U3647 : INV_X1 port map( A => n5846, ZN => n5847);
   U3648 : OAI21_X1 port map( B1 => n5847, B2 => n8423, A => n5879, ZN => n5851
                           );
   U3649 : NAND3_X1 port map( A1 => n367, A2 => n5848, A3 => n8423, ZN => n5849
                           );
   U3650 : NAND2_X1 port map( A1 => n8397, A2 => n5849, ZN => n5850);
   U3651 : NAND2_X1 port map( A1 => n5851, A2 => n5850, ZN => n5852);
   U3652 : NAND2_X1 port map( A1 => n5853, A2 => n5852, ZN => n6143);
   U3653 : MUX2_X1 port map( A => n6715, B => n6243, S => n360, Z => n5857);
   U3654 : XNOR2_X1 port map( A => n5854, B => n372, ZN => n5855);
   U3655 : NAND2_X1 port map( A1 => n7861, A2 => n5855, ZN => n5856);
   U3656 : NAND2_X1 port map( A1 => n5857, A2 => n5856, ZN => n6144);
   U3657 : XNOR2_X1 port map( A => n6143, B => n6144, ZN => n5860);
   U3658 : MUX2_X1 port map( A => n4490, B => n7051, S => n377, Z => n5859);
   U3659 : MUX2_X1 port map( A => n4607, B => n8595, S => n359, Z => n5858);
   U3660 : NAND2_X1 port map( A1 => n5859, A2 => n5858, ZN => n6140);
   U3661 : XNOR2_X1 port map( A => n5860, B => n6140, ZN => n6132);
   U3662 : XNOR2_X1 port map( A => n6132, B => n6136, ZN => n5871);
   U3663 : INV_X1 port map( A => n5861, ZN => n7047);
   U3664 : MUX2_X1 port map( A => n7047, B => n7665, S => n8401, Z => n5863);
   U3665 : MUX2_X1 port map( A => n7696, B => n7695, S => n8324, Z => n5862);
   U3666 : XNOR2_X1 port map( A => n8325, B => n8002, ZN => n5864);
   U3667 : INV_X1 port map( A => n5866, ZN => n7094);
   U3668 : INV_X1 port map( A => n5867, ZN => n7093);
   U3669 : MUX2_X1 port map( A => n7094, B => n7093, S => n362, Z => n5869);
   U3670 : INV_X1 port map( A => n6800, ZN => n7096);
   U3671 : INV_X1 port map( A => n6342, ZN => n7095);
   U3672 : NOR2_X1 port map( A1 => n5869, A2 => n5868, ZN => n6178);
   U3674 : XNOR2_X1 port map( A => n8498, B => n6174, ZN => n5870);
   U3675 : XNOR2_X1 port map( A => n5870, B => n6175, ZN => n6135);
   U3676 : INV_X1 port map( A => n6135, ZN => n6137);
   U3677 : MUX2_X1 port map( A => n5873, B => n5872, S => n377, Z => n5877);
   U3678 : XNOR2_X1 port map( A => n360, B => n6244, ZN => n5874);
   U3679 : NOR2_X1 port map( A1 => n5875, A2 => n5874, ZN => n5876);
   U3680 : NOR2_X1 port map( A1 => n5877, A2 => n5876, ZN => n5918);
   U3681 : MUX2_X1 port map( A => n6103, B => n6102, S => n8325, Z => n5882);
   U3682 : XNOR2_X1 port map( A => n5879, B => n8349, ZN => n5880);
   U3683 : NAND2_X1 port map( A1 => n5880, A2 => n6104, ZN => n5881);
   U3684 : NAND2_X1 port map( A1 => n5882, A2 => n5881, ZN => n5920);
   U3685 : MUX2_X1 port map( A => n8469, B => n8595, S => n356, Z => n5886);
   U3686 : XNOR2_X1 port map( A => n5883, B => n8394, ZN => n5884);
   U3687 : NAND2_X1 port map( A1 => n4491, A2 => n5884, ZN => n5885);
   U3688 : NAND2_X1 port map( A1 => n5886, A2 => n5885, ZN => n5887);
   U3689 : NAND2_X1 port map( A1 => n5920, A2 => n5887, ZN => n5889);
   U3691 : INV_X1 port map( A => n5887, ZN => n5921);
   U3693 : MUX2_X1 port map( A => n7121, B => n7120, S => n356, Z => n6187);
   U3694 : MUX2_X1 port map( A => n8593, B => n6812, S => n373, Z => n6183);
   U3695 : NAND2_X1 port map( A1 => n6187, A2 => n6183, ZN => n5891);
   U3696 : NAND2_X1 port map( A1 => n8504, A2 => n8393, ZN => n6184);
   U3697 : XNOR2_X1 port map( A => n6184, B => n6259, ZN => n5890);
   U3698 : XNOR2_X1 port map( A => n5891, B => n5890, ZN => n5892);
   U3699 : NAND2_X1 port map( A1 => n5893, A2 => n5892, ZN => n6201);
   U3700 : INV_X1 port map( A => n5892, ZN => n5895);
   U3702 : NAND2_X1 port map( A1 => n5895, A2 => n5894, ZN => n6202);
   U3703 : NAND2_X1 port map( A1 => n6201, A2 => n6202, ZN => n5908);
   U3704 : MUX2_X1 port map( A => n7053, B => n8501, S => n7945, Z => n5897);
   U3705 : MUX2_X1 port map( A => n4462, B => n7198, S => n8333, Z => n5896);
   U3706 : MUX2_X1 port map( A => n5898, B => n8535, S => n357, Z => n5900);
   U3707 : MUX2_X1 port map( A => n8454, B => n8515, S => n205, Z => n5899);
   U3708 : NAND2_X1 port map( A1 => n5900, A2 => n5899, ZN => n5903);
   U3709 : MUX2_X1 port map( A => n4487, B => n7325, S => n204, Z => n5902);
   U3710 : MUX2_X1 port map( A => n7324, B => n8465, S => B_SIG_9_port, Z => 
                           n5901);
   U3711 : NAND2_X1 port map( A1 => n5902, A2 => n5901, ZN => n5904);
   U3712 : NAND2_X1 port map( A1 => n5903, A2 => n5904, ZN => n5950);
   U3713 : NAND2_X1 port map( A1 => n5952, A2 => n5950, ZN => n5907);
   U3714 : INV_X1 port map( A => n5903, ZN => n5906);
   U3715 : INV_X1 port map( A => n5904, ZN => n5905);
   U3716 : NAND2_X1 port map( A1 => n5906, A2 => n5905, ZN => n5951);
   U3718 : XNOR2_X1 port map( A => n5908, B => n6199, ZN => n5909);
   U3719 : NAND2_X1 port map( A1 => n5910, A2 => n5909, ZN => n6212);
   U3720 : NAND2_X1 port map( A1 => n6212, A2 => n6211, ZN => n5933);
   U3721 : MUX2_X1 port map( A => n7086, B => n7047, S => n8324, Z => n5912);
   U3722 : MUX2_X1 port map( A => n8559, B => n7695, S => n386, Z => n5911);
   U3723 : NAND2_X1 port map( A1 => n5912, A2 => n5911, ZN => n5993);
   U3724 : INV_X1 port map( A => n6259, ZN => n6431);
   U3725 : NAND2_X1 port map( A1 => n6431, A2 => n7506, ZN => n5913);
   U3726 : AND2_X1 port map( A1 => n7947, A2 => n5913, ZN => n5990);
   U3727 : XNOR2_X1 port map( A => n5993, B => n5990, ZN => n5917);
   U3728 : MUX2_X1 port map( A => n8445, B => n6740, S => n363, Z => n5916);
   U3729 : MUX2_X1 port map( A => n8459, B => n8434, S => n8330, Z => n5915);
   U3730 : NAND2_X1 port map( A1 => n5916, A2 => n5915, ZN => n5991);
   U3731 : XNOR2_X1 port map( A => n5917, B => n5991, ZN => n5928);
   U3732 : INV_X1 port map( A => n5918, ZN => n5919);
   U3733 : XNOR2_X1 port map( A => n5920, B => n5919, ZN => n5922);
   U3734 : XNOR2_X1 port map( A => n5922, B => n5921, ZN => n5929);
   U3735 : NAND2_X1 port map( A1 => n5928, A2 => n5929, ZN => n5964);
   U3736 : INV_X1 port map( A => n5923, ZN => n5925);
   U3737 : NAND2_X1 port map( A1 => n5925, A2 => n5924, ZN => n5927);
   U3738 : NAND2_X1 port map( A1 => n5927, A2 => n5926, ZN => n5966);
   U3739 : NAND2_X1 port map( A1 => n5964, A2 => n5966, ZN => n5932);
   U3740 : INV_X1 port map( A => n5928, ZN => n5931);
   U3741 : INV_X1 port map( A => n5929, ZN => n5930);
   U3742 : NAND2_X1 port map( A1 => n5931, A2 => n5930, ZN => n5965);
   U3743 : NAND2_X1 port map( A1 => n5932, A2 => n5965, ZN => n6210);
   U3744 : XNOR2_X1 port map( A => n5933, B => n6210, ZN => n6218);
   U3745 : AND2_X1 port map( A1 => n5935, A2 => n5934, ZN => n5997);
   U3746 : NAND2_X2 port map( A1 => n5937, A2 => n5936, ZN => n7253);
   U3748 : MUX2_X1 port map( A => n7253, B => n7771, S => n381, Z => n5939);
   U3749 : MUX2_X1 port map( A => n7692, B => n7773, S => n8393, Z => n5938);
   U3750 : NAND2_X1 port map( A1 => n5939, A2 => n5938, ZN => n5996);
   U3751 : XNOR2_X1 port map( A => n5997, B => n5996, ZN => n5949);
   U3752 : INV_X1 port map( A => n5947, ZN => n5944);
   U3753 : INV_X1 port map( A => n5940, ZN => n5942);
   U3754 : AOI21_X1 port map( B1 => n5942, B2 => n5947, A => n5941, ZN => n5943
                           );
   U3755 : OAI21_X1 port map( B1 => n5945, B2 => n5944, A => n5943, ZN => n5946
                           );
   U3756 : OAI21_X1 port map( B1 => n5948, B2 => n5947, A => n5946, ZN => n5998
                           );
   U3757 : XNOR2_X1 port map( A => n5949, B => n5998, ZN => n5954);
   U3758 : NAND2_X1 port map( A1 => n5951, A2 => n5950, ZN => n5953);
   U3759 : XNOR2_X1 port map( A => n5953, B => n5952, ZN => n5955);
   U3760 : NAND2_X1 port map( A1 => n5954, A2 => n5955, ZN => n6031);
   U3761 : INV_X1 port map( A => n5954, ZN => n5956);
   U3762 : NAND2_X1 port map( A1 => n5956, A2 => n4497, ZN => n6029);
   U3763 : NAND2_X1 port map( A1 => n6031, A2 => n6029, ZN => n5963);
   U3764 : INV_X1 port map( A => n5957, ZN => n5962);
   U3765 : INV_X1 port map( A => n5958, ZN => n5961);
   U3766 : INV_X1 port map( A => n5959, ZN => n5960);
   U3767 : FA_X1 port map( A => n5962, B => n5961, CI => n5960, CO => n6028, S 
                           => n_1138);
   U3768 : XNOR2_X1 port map( A => n8557, B => n8531, ZN => n5978);
   U3769 : NAND2_X1 port map( A1 => n5965, A2 => n5964, ZN => n5967);
   U3770 : XNOR2_X1 port map( A => n5967, B => n5966, ZN => n5979);
   U3771 : NAND2_X1 port map( A1 => n5978, A2 => n5979, ZN => n6059);
   U3772 : INV_X1 port map( A => n5968, ZN => n5969);
   U3773 : NAND2_X1 port map( A1 => n5732, A2 => n5969, ZN => n5974);
   U3774 : INV_X1 port map( A => n5971, ZN => n5977);
   U3775 : INV_X1 port map( A => n5970, ZN => n5973);
   U3776 : NAND2_X1 port map( A1 => n5971, A2 => n5973, ZN => n5976);
   U3777 : NAND3_X1 port map( A1 => n5974, A2 => n5973, A3 => n5972, ZN => 
                           n5975);
   U3778 : NAND2_X1 port map( A1 => n6059, A2 => n6076, ZN => n5981);
   U3779 : INV_X1 port map( A => n5979, ZN => n5980);
   U3780 : NAND2_X1 port map( A1 => n4496, A2 => n5980, ZN => n6060);
   U3781 : NAND2_X1 port map( A1 => n5981, A2 => n6060, ZN => n6217);
   U3782 : XNOR2_X1 port map( A => n6218, B => n6217, ZN => n6053);
   U3783 : MUX2_X1 port map( A => n7121, B => n4360, S => n373, Z => n5983);
   U3784 : MUX2_X1 port map( A => n8593, B => n7122, S => n379, Z => n5982);
   U3785 : NAND2_X1 port map( A1 => n5983, A2 => n5982, ZN => n6008);
   U3787 : AND2_X1 port map( A1 => A_SIG_23_port, A2 => n8354, ZN => n6005);
   U3788 : MUX2_X1 port map( A => n8476, B => n7559, S => n390, Z => n5985);
   U3789 : MUX2_X1 port map( A => n7227, B => n7439, S => n6606, Z => n5984);
   U3790 : NAND2_X1 port map( A1 => n5985, A2 => n5984, ZN => n6007);
   U3791 : OAI21_X1 port map( B1 => n6008, B2 => n6005, A => n6007, ZN => n5987
                           );
   U3792 : NAND2_X1 port map( A1 => n6008, A2 => n6005, ZN => n5986);
   U3793 : NAND2_X1 port map( A1 => n5987, A2 => n5986, ZN => n6163);
   U3794 : MUX2_X1 port map( A => n7253, B => n7392, S => n386, Z => n5989);
   U3795 : MUX2_X1 port map( A => n7692, B => n7773, S => n8396, Z => n5988);
   U3797 : XNOR2_X1 port map( A => n6163, B => n6171, ZN => n5995);
   U3798 : INV_X1 port map( A => n5990, ZN => n5992);
   U3799 : NOR2_X1 port map( A1 => n5993, A2 => n5992, ZN => n6165);
   U3800 : INV_X1 port map( A => n5991, ZN => n5994);
   U3801 : NAND2_X1 port map( A1 => n5993, A2 => n5992, ZN => n6164);
   U3802 : XNOR2_X1 port map( A => n6162, B => n5995, ZN => n6001);
   U3803 : INV_X1 port map( A => n5996, ZN => n6000);
   U3804 : INV_X1 port map( A => n5997, ZN => n5999);
   U3805 : FA_X1 port map( A => n6000, B => n5999, CI => n5998, CO => n6002, S 
                           => n_1139);
   U3806 : NAND2_X1 port map( A1 => n6001, A2 => n6002, ZN => n6208);
   U3807 : INV_X1 port map( A => n6001, ZN => n6004);
   U3808 : INV_X1 port map( A => n6002, ZN => n6003);
   U3809 : NAND2_X1 port map( A1 => n6004, A2 => n6003, ZN => n6207);
   U3810 : NAND2_X1 port map( A1 => n6208, A2 => n6207, ZN => n6027);
   U3811 : INV_X1 port map( A => n6005, ZN => n6006);
   U3812 : XNOR2_X1 port map( A => n6007, B => n6006, ZN => n6010);
   U3813 : INV_X1 port map( A => n6008, ZN => n6009);
   U3814 : XNOR2_X1 port map( A => n6010, B => n6009, ZN => n6022);
   U3815 : INV_X1 port map( A => n6011, ZN => n6014);
   U3816 : AOI21_X1 port map( B1 => n6014, B2 => n6013, A => n6012, ZN => n6016
                           );
   U3817 : NOR2_X1 port map( A1 => n6014, A2 => n6013, ZN => n6015);
   U3818 : NOR2_X1 port map( A1 => n6016, A2 => n6015, ZN => n6023);
   U3819 : NAND2_X1 port map( A1 => n6022, A2 => n6023, ZN => n6033);
   U3820 : INV_X1 port map( A => n6017, ZN => n6018);
   U3821 : NAND2_X1 port map( A1 => n6019, A2 => n6018, ZN => n6021);
   U3822 : NAND2_X1 port map( A1 => n6021, A2 => n6020, ZN => n6035);
   U3823 : NAND2_X1 port map( A1 => n6033, A2 => n6035, ZN => n6026);
   U3824 : INV_X1 port map( A => n6022, ZN => n6025);
   U3825 : INV_X1 port map( A => n6023, ZN => n6024);
   U3826 : NAND2_X1 port map( A1 => n6025, A2 => n6024, ZN => n6034);
   U3827 : NAND2_X1 port map( A1 => n6026, A2 => n6034, ZN => n6206);
   U3828 : INV_X1 port map( A => n6028, ZN => n6030);
   U3829 : NAND2_X1 port map( A1 => n6030, A2 => n6029, ZN => n6032);
   U3831 : XNOR2_X1 port map( A => n6522, B => n6521, ZN => n6052);
   U3832 : NAND2_X1 port map( A1 => n6034, A2 => n6033, ZN => n6037);
   U3833 : INV_X1 port map( A => n6035, ZN => n6036);
   U3834 : XNOR2_X1 port map( A => n6037, B => n6036, ZN => n6049);
   U3835 : INV_X1 port map( A => n6038, ZN => n6042);
   U3836 : NAND2_X1 port map( A1 => n6046, A2 => n6045, ZN => n6048);
   U3837 : NAND2_X1 port map( A1 => n6048, A2 => n6047, ZN => n6058);
   U3838 : NAND2_X1 port map( A1 => n6057, A2 => n6058, ZN => n6093);
   U3839 : INV_X1 port map( A => n6050, ZN => n6051);
   U3840 : NAND2_X1 port map( A1 => n4434, A2 => n6051, ZN => n6091);
   U3842 : XNOR2_X1 port map( A => n6221, B => n6053, ZN => n8049);
   U3843 : NAND2_X1 port map( A1 => n6091, A2 => n6057, ZN => n6080);
   U3844 : INV_X1 port map( A => n6058, ZN => n6075);
   U3845 : XNOR2_X1 port map( A => n6080, B => n6075, ZN => n6063);
   U3846 : NAND2_X1 port map( A1 => n6060, A2 => n6059, ZN => n6081);
   U3847 : INV_X1 port map( A => n6076, ZN => n6061);
   U3848 : XNOR2_X1 port map( A => n6081, B => n6061, ZN => n6062);
   U3849 : NAND2_X1 port map( A1 => n8049, A2 => n8050, ZN => n8048);
   U3850 : INV_X1 port map( A => n6064, ZN => n6066);
   U3851 : NAND2_X1 port map( A1 => n6066, A2 => n4464, ZN => n8032);
   U3852 : INV_X1 port map( A => n6073, ZN => n6067);
   U3853 : NAND2_X1 port map( A1 => n6067, A2 => n6068, ZN => n6070);
   U3854 : INV_X1 port map( A => n6068, ZN => n6069);
   U3855 : AOI22_X1 port map( A1 => n6074, A2 => n6070, B1 => n6069, B2 => 
                           n6073, ZN => n8040);
   U3856 : INV_X1 port map( A => n6071, ZN => n6072);
   U3857 : OAI21_X1 port map( B1 => n6074, B2 => n6073, A => n6072, ZN => n8042
                           );
   U3859 : XNOR2_X1 port map( A => n6076, B => n6075, ZN => n6079);
   U3860 : INV_X1 port map( A => n6077, ZN => n6078);
   U3861 : XNOR2_X1 port map( A => n6079, B => n6078, ZN => n6083);
   U3862 : XNOR2_X1 port map( A => n8532, B => n6080, ZN => n6082);
   U3864 : NAND2_X1 port map( A1 => n7943, A2 => n7940, ZN => n6084);
   U3866 : OAI21_X1 port map( B1 => n7940, B2 => n7943, A => n8050, ZN => n6090
                           );
   U3867 : INV_X1 port map( A => n8049, ZN => n6089);
   U3868 : AND2_X1 port map( A1 => n6090, A2 => n6089, ZN => n7619);
   U3869 : NOR3_X1 port map( A1 => n8050, A2 => n7943, A3 => n7940, ZN => n7620
                           );
   U3871 : NAND2_X1 port map( A1 => n8204, A2 => n8209, ZN => n8121);
   U3872 : NAND2_X1 port map( A1 => n4433, A2 => n6521, ZN => n6096);
   U3873 : INV_X1 port map( A => n6521, ZN => n6092);
   U3874 : NAND3_X1 port map( A1 => n6093, A2 => n6092, A3 => n6091, ZN => 
                           n6094);
   U3875 : NAND2_X1 port map( A1 => n6094, A2 => n6522, ZN => n6095);
   U3876 : MUX2_X1 port map( A => n4489, B => n7084, S => n360, Z => n6098);
   U3877 : MUX2_X1 port map( A => n8469, B => n8596, S => n377, Z => n6097);
   U3878 : NAND2_X1 port map( A1 => n6098, A2 => n6097, ZN => n6281);
   U3879 : MUX2_X1 port map( A => n6715, B => n6243, S => n372, Z => n6101);
   U3880 : XNOR2_X1 port map( A => n8329, B => n6244, ZN => n6099);
   U3881 : NAND2_X1 port map( A1 => n7861, A2 => n6099, ZN => n6100);
   U3882 : NAND2_X1 port map( A1 => n6101, A2 => n6100, ZN => n6280);
   U3883 : MUX2_X1 port map( A => n6103, B => n6102, S => n8334, Z => n6107);
   U3884 : XNOR2_X1 port map( A => n4809, B => n357, ZN => n6252);
   U3885 : INV_X1 port map( A => n6252, ZN => n6105);
   U3886 : NAND2_X1 port map( A1 => n6105, A2 => n6104, ZN => n6106);
   U3887 : NAND2_X1 port map( A1 => n6107, A2 => n6106, ZN => n6279);
   U3888 : MUX2_X1 port map( A => n6800, B => n6342, S => n362, Z => n6112);
   U3889 : XNOR2_X1 port map( A => n6109, B => n6593, ZN => n6110);
   U3890 : NAND2_X1 port map( A1 => n6110, A2 => n6595, ZN => n6111);
   U3891 : MUX2_X1 port map( A => n8559, B => n8582, S => n6606, Z => n6117);
   U3892 : XNOR2_X1 port map( A => n6234, B => n390, ZN => n6114);
   U3893 : NAND2_X1 port map( A1 => n6374, A2 => n6114, ZN => n6116);
   U3894 : AND2_X1 port map( A1 => n6117, A2 => n6116, ZN => n6119);
   U3895 : NAND2_X1 port map( A1 => n6118, A2 => n6119, ZN => n6299);
   U3896 : INV_X1 port map( A => n6119, ZN => n6120);
   U3897 : NAND2_X1 port map( A1 => n6121, A2 => n6120, ZN => n6296);
   U3898 : NAND2_X1 port map( A1 => n6299, A2 => n6296, ZN => n6123);
   U3899 : MUX2_X1 port map( A => n8445, B => n6740, S => n8423, Z => n6298);
   U3900 : MUX2_X1 port map( A => n8459, B => n8434, S => n8325, Z => n6297);
   U3901 : NAND2_X1 port map( A1 => n6298, A2 => n6297, ZN => n6122);
   U3902 : XNOR2_X1 port map( A => n6123, B => n6122, ZN => n6267);
   U3903 : XNOR2_X1 port map( A => n6268, B => n6267, ZN => n6131);
   U3904 : MUX2_X1 port map( A => n7324, B => n8465, S => n8392, Z => n6124);
   U3905 : NAND2_X1 port map( A1 => n6125, A2 => n6124, ZN => n6283);
   U3906 : MUX2_X1 port map( A => n8454, B => n8516, S => n7506, Z => n6127);
   U3908 : XNOR2_X1 port map( A => n6283, B => n6284, ZN => n6130);
   U3909 : MUX2_X1 port map( A => n8500, B => n7053, S => n204, Z => n6129);
   U3910 : MUX2_X1 port map( A => n4462, B => n7054, S => B_SIG_9_port, Z => 
                           n6128);
   U3911 : NAND2_X1 port map( A1 => n6129, A2 => n6128, ZN => n6285);
   U3912 : XNOR2_X1 port map( A => n6285, B => n6130, ZN => n6269);
   U3913 : XNOR2_X1 port map( A => n6131, B => n6269, ZN => n6504);
   U3915 : INV_X1 port map( A => n6132, ZN => n6133);
   U3916 : OAI21_X1 port map( B1 => n6135, B2 => n8572, A => n6133, ZN => n6139
                           );
   U3917 : OR2_X1 port map( A1 => n6137, A2 => n6136, ZN => n6138);
   U3918 : NAND2_X1 port map( A1 => n6138, A2 => n6139, ZN => n6506);
   U3919 : INV_X1 port map( A => n6140, ZN => n6142);
   U3920 : NAND2_X1 port map( A1 => n6143, A2 => n6144, ZN => n6141);
   U3921 : NAND2_X1 port map( A1 => n6142, A2 => n6141, ZN => n6148);
   U3922 : INV_X1 port map( A => n6143, ZN => n6146);
   U3923 : INV_X1 port map( A => n6144, ZN => n6145);
   U3924 : NAND2_X1 port map( A1 => n6146, A2 => n6145, ZN => n6147);
   U3925 : NAND2_X1 port map( A1 => n6148, A2 => n6147, ZN => n6324);
   U3926 : INV_X1 port map( A => n6149, ZN => n6151);
   U3927 : INV_X1 port map( A => n6152, ZN => n6155);
   U3928 : INV_X1 port map( A => n6153, ZN => n6154);
   U3929 : NAND2_X1 port map( A1 => n6155, A2 => n6154, ZN => n6156);
   U3930 : NAND2_X1 port map( A1 => n6157, A2 => n6156, ZN => n6325);
   U3931 : XNOR2_X1 port map( A => n6325, B => n6324, ZN => n6160);
   U3932 : MUX2_X1 port map( A => n8593, B => n6812, S => n356, Z => n6303);
   U3933 : NAND2_X1 port map( A1 => n6307, A2 => n6303, ZN => n6159);
   U3934 : AND2_X1 port map( A1 => n8504, A2 => n8396, ZN => n6301);
   U3935 : INV_X1 port map( A => n6301, ZN => n6304);
   U3936 : XNOR2_X1 port map( A => n6304, B => n6431, ZN => n6158);
   U3937 : XNOR2_X1 port map( A => n6159, B => n6158, ZN => n6326);
   U3938 : XNOR2_X1 port map( A => n6160, B => n6326, ZN => n6503);
   U3939 : INV_X1 port map( A => n6503, ZN => n6507);
   U3940 : XNOR2_X1 port map( A => n6506, B => n6507, ZN => n6161);
   U3941 : XNOR2_X1 port map( A => n6504, B => n6161, ZN => n6524);
   U3942 : INV_X1 port map( A => n6163, ZN => n6170);
   U3943 : INV_X1 port map( A => n6164, ZN => n6168);
   U3944 : INV_X1 port map( A => n6165, ZN => n6167);
   U3945 : INV_X1 port map( A => n6171, ZN => n6166);
   U3946 : OAI211_X1 port map( C1 => n6168, C2 => n5991, A => n6167, B => n6166
                           , ZN => n6169);
   U3947 : AOI22_X1 port map( A1 => n6172, A2 => n6171, B1 => n6169, B2 => 
                           n6170, ZN => n6196);
   U3948 : NAND2_X1 port map( A1 => n6174, A2 => n8498, ZN => n6176);
   U3949 : NAND2_X1 port map( A1 => n6176, A2 => n6175, ZN => n6180);
   U3950 : NAND2_X1 port map( A1 => n6178, A2 => n6177, ZN => n6179);
   U3951 : NAND2_X1 port map( A1 => n6180, A2 => n6179, ZN => n6334);
   U3952 : INV_X1 port map( A => n6334, ZN => n6195);
   U3953 : INV_X1 port map( A => n6184, ZN => n6181);
   U3954 : NAND2_X1 port map( A1 => n6181, A2 => n6431, ZN => n6182);
   U3955 : AND2_X1 port map( A1 => n6183, A2 => n6182, ZN => n6186);
   U3956 : AND2_X1 port map( A1 => n6184, A2 => n6259, ZN => n6185);
   U3957 : AOI21_X1 port map( B1 => n6186, B2 => n6187, A => n6185, ZN => n6193
                           );
   U3958 : INV_X1 port map( A => n6193, ZN => n6191);
   U3959 : MUX2_X1 port map( A => n7253, B => n7392, S => n8324, Z => n6189);
   U3960 : MUX2_X1 port map( A => n7692, B => n7773, S => n8328, Z => n6188);
   U3961 : NAND2_X1 port map( A1 => n6189, A2 => n6188, ZN => n6192);
   U3962 : INV_X1 port map( A => n6192, ZN => n6190);
   U3963 : NAND2_X1 port map( A1 => n6191, A2 => n6190, ZN => n6335);
   U3964 : NAND2_X1 port map( A1 => n6193, A2 => n6192, ZN => n6333);
   U3965 : NAND2_X1 port map( A1 => n6335, A2 => n6333, ZN => n6194);
   U3966 : XNOR2_X1 port map( A => n6195, B => n6194, ZN => n6197);
   U3967 : NAND2_X1 port map( A1 => n6197, A2 => n8591, ZN => n6501);
   U3968 : NOR2_X1 port map( A1 => n6197, A2 => n6196, ZN => n6499);
   U3969 : INV_X1 port map( A => n6499, ZN => n6198);
   U3970 : NAND2_X1 port map( A1 => n6198, A2 => n6501, ZN => n6205);
   U3971 : INV_X1 port map( A => n6199, ZN => n6200);
   U3972 : NAND2_X1 port map( A1 => n6201, A2 => n6200, ZN => n6203);
   U3973 : NAND2_X1 port map( A1 => n6203, A2 => n6202, ZN => n6500);
   U3974 : INV_X1 port map( A => n6500, ZN => n6204);
   U3975 : XNOR2_X1 port map( A => n6205, B => n6204, ZN => n6516);
   U3976 : NAND2_X1 port map( A1 => n6207, A2 => n6206, ZN => n6209);
   U3977 : NAND2_X1 port map( A1 => n6209, A2 => n6208, ZN => n6539);
   U3978 : XNOR2_X1 port map( A => n6516, B => n6539, ZN => n6215);
   U3979 : NAND2_X1 port map( A1 => n6211, A2 => n6210, ZN => n6213);
   U3980 : NAND2_X1 port map( A1 => n6213, A2 => n6212, ZN => n6517);
   U3981 : XNOR2_X1 port map( A => n6215, B => n6214, ZN => n6525);
   U3982 : INV_X1 port map( A => n6217, ZN => n6219);
   U3984 : NAND2_X1 port map( A1 => n6223, A2 => n6224, ZN => n8073);
   U3985 : MUX2_X1 port map( A => n4490, B => n8577, S => n372, Z => n6226);
   U3986 : MUX2_X1 port map( A => n8469, B => n8596, S => n360, Z => n6225);
   U3987 : NAND2_X1 port map( A1 => n6226, A2 => n6225, ZN => n6440);
   U3988 : INV_X1 port map( A => n6227, ZN => n6228);
   U3989 : OAI21_X1 port map( B1 => n6228, B2 => n204, A => n6706, ZN => n6233)
                           ;
   U3990 : NAND3_X1 port map( A1 => n8353, A2 => n6229, A3 => n204, ZN => n6230
                           );
   U3991 : NAND2_X1 port map( A1 => n6230, A2 => n8357, ZN => n6232);
   U3992 : XNOR2_X1 port map( A => n8392, B => n6705, ZN => n6231);
   U3993 : AOI22_X1 port map( A1 => n6233, A2 => n6232, B1 => n6231, B2 => 
                           n6702, ZN => n6238);
   U3994 : NAND2_X1 port map( A1 => n8582, A2 => n390, ZN => n6237);
   U3995 : NAND2_X1 port map( A1 => n8559, A2 => n8352, ZN => n6236);
   U3996 : XNOR2_X1 port map( A => n6234, B => n362, ZN => n6235);
   U3997 : AOI22_X1 port map( A1 => n6237, A2 => n6236, B1 => n6374, B2 => 
                           n6235, ZN => n6239);
   U3998 : NAND2_X1 port map( A1 => n6238, A2 => n6239, ZN => n6438);
   U4002 : NAND2_X1 port map( A1 => n6438, A2 => n6437, ZN => n6242);
   U4004 : MUX2_X1 port map( A => n6715, B => n6243, S => n363, Z => n6247);
   U4005 : XNOR2_X1 port map( A => n8325, B => n6244, ZN => n6245);
   U4006 : NAND2_X1 port map( A1 => n7861, A2 => n6245, ZN => n6246);
   U4007 : NAND2_X1 port map( A1 => n6247, A2 => n6246, ZN => n6424);
   U4008 : NAND2_X1 port map( A1 => n6249, A2 => n8516, ZN => n6427);
   U4009 : XNOR2_X1 port map( A => n5879, B => n8363, ZN => n6250);
   U4010 : NAND2_X1 port map( A1 => n6250, A2 => n6251, ZN => n6381);
   U4011 : XNOR2_X1 port map( A => n5879, B => n7769, ZN => n6382);
   U4013 : XNOR2_X1 port map( A => n6427, B => n8429, ZN => n6253);
   U4014 : XNOR2_X1 port map( A => n6253, B => n6424, ZN => n6442);
   U4015 : XNOR2_X1 port map( A => n6445, B => n6442, ZN => n6266);
   U4016 : NAND2_X1 port map( A1 => n6688, A2 => n4381, ZN => n6255);
   U4017 : NAND2_X1 port map( A1 => n7324, A2 => n373, ZN => n6254);
   U4018 : NAND2_X1 port map( A1 => n6255, A2 => n6254, ZN => n6258);
   U4019 : XNOR2_X1 port map( A => n8326, B => n6229, ZN => n6256);
   U4020 : NAND2_X1 port map( A1 => n5041, A2 => n6256, ZN => n6257);
   U4021 : NAND2_X1 port map( A1 => n6258, A2 => n6257, ZN => n6430);
   U4022 : XNOR2_X1 port map( A => n6430, B => n6259, ZN => n6265);
   U4023 : XNOR2_X1 port map( A => n8334, B => n8002, ZN => n6263);
   U4024 : OAI21_X1 port map( B1 => n6743, B2 => n8349, A => n4809, ZN => n6262
                           );
   U4025 : NAND3_X1 port map( A1 => n8335, A2 => n8349, A3 => n8002, ZN => 
                           n6260);
   U4026 : NAND2_X1 port map( A1 => n8397, A2 => n6260, ZN => n6261);
   U4027 : AOI22_X1 port map( A1 => n6264, A2 => n6263, B1 => n6262, B2 => 
                           n6261, ZN => n6434);
   U4028 : XNOR2_X1 port map( A => n6265, B => n6434, ZN => n6443);
   U4029 : OAI21_X1 port map( B1 => n6269, B2 => n6268, A => n6267, ZN => n6271
                           );
   U4030 : NAND2_X1 port map( A1 => n6269, A2 => n6268, ZN => n6270);
   U4031 : NAND2_X1 port map( A1 => n6271, A2 => n6270, ZN => n6534);
   U4032 : MUX2_X1 port map( A => n6342, B => n6800, S => n6109, Z => n6274);
   U4033 : XNOR2_X1 port map( A => B_SIG_9_port, B => n6343, ZN => n6272);
   U4034 : NAND2_X1 port map( A1 => n6272, A2 => n6595, ZN => n6273);
   U4035 : NAND2_X1 port map( A1 => n6273, A2 => n6274, ZN => n6318);
   U4036 : NAND2_X1 port map( A1 => n4514, A2 => n8328, ZN => n6317);
   U4037 : XNOR2_X1 port map( A => n6318, B => n6317, ZN => n6278);
   U4038 : MUX2_X1 port map( A => n7121, B => n4360, S => n377, Z => n6277);
   U4039 : MUX2_X1 port map( A => n8593, B => n7122, S => n359, Z => n6276);
   U4040 : NAND2_X1 port map( A1 => n6277, A2 => n6276, ZN => n6320);
   U4041 : XNOR2_X1 port map( A => n6278, B => n6320, ZN => n6293);
   U4042 : AND2_X1 port map( A1 => n6279, A2 => n6280, ZN => n6282);
   U4043 : OAI22_X1 port map( A1 => n6282, A2 => n6281, B1 => n6280, B2 => 
                           n6279, ZN => n6291);
   U4044 : XNOR2_X1 port map( A => n6293, B => n6291, ZN => n6288);
   U4045 : OAI21_X1 port map( B1 => n6285, B2 => n6284, A => n6283, ZN => n6287
                           );
   U4046 : NAND2_X1 port map( A1 => n6285, A2 => n6284, ZN => n6286);
   U4048 : NAND2_X1 port map( A1 => n6293, A2 => n6292, ZN => n6294);
   U4049 : NAND2_X1 port map( A1 => n6295, A2 => n6294, ZN => n6454);
   U4050 : NAND3_X1 port map( A1 => n6298, A2 => n6297, A3 => n6296, ZN => 
                           n6300);
   U4051 : NAND2_X1 port map( A1 => n6300, A2 => n6299, ZN => n6331);
   U4052 : NAND2_X1 port map( A1 => n6301, A2 => n6431, ZN => n6302);
   U4053 : AND2_X1 port map( A1 => n6303, A2 => n6302, ZN => n6306);
   U4054 : AND2_X1 port map( A1 => n6304, A2 => n6259, ZN => n6305);
   U4056 : MUX2_X1 port map( A => n7253, B => n7392, S => n376, Z => n6309);
   U4057 : MUX2_X1 port map( A => n7692, B => n7773, S => n8350, Z => n6308);
   U4058 : NAND2_X1 port map( A1 => n6309, A2 => n6308, ZN => n6311);
   U4059 : NAND2_X1 port map( A1 => n6310, A2 => n6311, ZN => n6329);
   U4060 : NAND2_X1 port map( A1 => n6331, A2 => n6329, ZN => n6312);
   U4061 : NAND2_X1 port map( A1 => n6312, A2 => n6330, ZN => n6452);
   U4062 : XNOR2_X1 port map( A => n6454, B => n6452, ZN => n6323);
   U4063 : MUX2_X1 port map( A => n6714, B => n6888, S => n8423, Z => n6314);
   U4064 : MUX2_X1 port map( A => n6715, B => n6887, S => n371, Z => n6313);
   U4065 : NAND2_X1 port map( A1 => n6314, A2 => n6313, ZN => n6477);
   U4066 : MUX2_X1 port map( A => n7253, B => n7771, S => n390, Z => n6316);
   U4067 : MUX2_X1 port map( A => n7692, B => n7773, S => n8401, Z => n6315);
   U4068 : NAND2_X1 port map( A1 => n6316, A2 => n6315, ZN => n6476);
   U4069 : XNOR2_X1 port map( A => n6477, B => n6476, ZN => n6322);
   U4070 : INV_X1 port map( A => n6317, ZN => n6319);
   U4071 : OAI21_X1 port map( B1 => n6320, B2 => n6319, A => n6318, ZN => n6475
                           );
   U4072 : NAND2_X1 port map( A1 => n6320, A2 => n6319, ZN => n6474);
   U4073 : NAND2_X1 port map( A1 => n6475, A2 => n6474, ZN => n6321);
   U4074 : XNOR2_X1 port map( A => n6322, B => n6321, ZN => n6451);
   U4075 : XNOR2_X1 port map( A => n6323, B => n6451, ZN => n6547);
   U4076 : NAND2_X1 port map( A1 => n6544, A2 => n6547, ZN => n6489);
   U4077 : OAI21_X1 port map( B1 => n6325, B2 => n6326, A => n6324, ZN => n6328
                           );
   U4078 : NAND2_X1 port map( A1 => n6326, A2 => n6325, ZN => n6327);
   U4079 : NAND2_X1 port map( A1 => n6328, A2 => n6327, ZN => n6496);
   U4080 : NAND2_X1 port map( A1 => n6332, A2 => n6338, ZN => n6337);
   U4081 : NAND2_X1 port map( A1 => n6334, A2 => n6333, ZN => n6336);
   U4082 : NAND2_X1 port map( A1 => n6336, A2 => n6335, ZN => n6495);
   U4083 : NAND2_X1 port map( A1 => n6337, A2 => n6495, ZN => n6340);
   U4084 : INV_X1 port map( A => n6338, ZN => n6497);
   U4085 : NAND2_X1 port map( A1 => n6497, A2 => n6496, ZN => n6339);
   U4086 : NAND2_X1 port map( A1 => n6489, A2 => n6548, ZN => n6341);
   U4087 : NAND2_X1 port map( A1 => n6341, A2 => n6490, ZN => n6668);
   U4088 : MUX2_X1 port map( A => n6800, B => n6342, S => n204, Z => n6346);
   U4089 : XNOR2_X1 port map( A => n6343, B => n8392, ZN => n6344);
   U4090 : NAND2_X1 port map( A1 => n6595, A2 => n6344, ZN => n6345);
   U4091 : AND2_X1 port map( A1 => n6346, A2 => n6345, ZN => n6350);
   U4092 : MUX2_X1 port map( A => n8582, B => n7090, S => B_SIG_8_port, Z => 
                           n6349);
   U4093 : XNOR2_X1 port map( A => B_SIG_9_port, B => n8503, ZN => n6347);
   U4094 : NAND2_X1 port map( A1 => n6374, A2 => n6347, ZN => n6348);
   U4095 : AND2_X1 port map( A1 => n6348, A2 => n6349, ZN => n6351);
   U4096 : NAND2_X1 port map( A1 => n6350, A2 => n6351, ZN => n6621);
   U4097 : NAND2_X1 port map( A1 => n6620, A2 => n6621, ZN => n6353);
   U4098 : MUX2_X1 port map( A => n8445, B => n6740, S => n7506, Z => n6619);
   U4099 : MUX2_X1 port map( A => n8459, B => n8434, S => n8331, Z => n6618);
   U4100 : NAND2_X1 port map( A1 => n6619, A2 => n6618, ZN => n6352);
   U4101 : XNOR2_X1 port map( A => n6353, B => n6352, ZN => n6602);
   U4102 : MUX2_X1 port map( A => n6811, B => n7120, S => n372, Z => n6605);
   U4103 : NAND2_X1 port map( A1 => n6605, A2 => n6608, ZN => n6356);
   U4104 : NAND2_X1 port map( A1 => n8504, A2 => n8350, ZN => n6409);
   U4105 : NAND2_X1 port map( A1 => n4514, A2 => n8401, ZN => n6354);
   U4106 : XNOR2_X1 port map( A => n6409, B => n6354, ZN => n6355);
   U4107 : XNOR2_X1 port map( A => n6356, B => n6355, ZN => n6948);
   U4108 : XNOR2_X1 port map( A => n6602, B => n6948, ZN => n6360);
   U4109 : MUX2_X1 port map( A => n8500, B => n7053, S => n356, Z => n6358);
   U4110 : MUX2_X1 port map( A => n4461, B => n7054, S => n4381, Z => n6357);
   U4111 : INV_X1 port map( A => n6591, ZN => n6589);
   U4112 : XNOR2_X1 port map( A => n6587, B => n6589, ZN => n6359);
   U4113 : MUX2_X1 port map( A => n4490, B => n8577, S => n371, Z => n6588);
   U4114 : MUX2_X1 port map( A => n8469, B => n8596, S => n363, Z => n6590);
   U4115 : XNOR2_X1 port map( A => n6359, B => n6592, ZN => n6949);
   U4116 : XNOR2_X1 port map( A => n6949, B => n6360, ZN => n6664);
   U4118 : XNOR2_X1 port map( A => n373, B => n6363, ZN => n6364);
   U4119 : NOR2_X1 port map( A1 => n6365, A2 => n6364, ZN => n6366);
   U4120 : MUX2_X1 port map( A => n8469, B => n8595, S => n372, Z => n6398);
   U4121 : XNOR2_X1 port map( A => n5883, B => n8329, ZN => n6368);
   U4122 : NAND2_X1 port map( A1 => n4491, A2 => n6368, ZN => n6396);
   U4123 : AND2_X1 port map( A1 => n6398, A2 => n6396, ZN => n6394);
   U4124 : XNOR2_X1 port map( A => n6395, B => n8470, ZN => n6370);
   U4125 : MUX2_X1 port map( A => n7324, B => n8465, S => n8326, Z => n6397);
   U4126 : NAND2_X1 port map( A1 => n6399, A2 => n6397, ZN => n6403);
   U4127 : INV_X1 port map( A => n6403, ZN => n6369);
   U4128 : XNOR2_X1 port map( A => n6370, B => n6369, ZN => n6420);
   U4129 : MUX2_X1 port map( A => n6800, B => n6342, S => n8327, Z => n6373);
   U4130 : XNOR2_X1 port map( A => n8351, B => n6593, ZN => n6371);
   U4131 : NAND2_X1 port map( A1 => n6595, A2 => n6371, ZN => n6372);
   U4132 : NAND2_X1 port map( A1 => n6373, A2 => n6372, ZN => n6380);
   U4133 : MUX2_X1 port map( A => n8559, B => n8582, S => n362, Z => n6377);
   U4134 : XNOR2_X1 port map( A => B_SIG_8_port, B => n5777, ZN => n6375);
   U4135 : NAND2_X1 port map( A1 => n6375, A2 => n6374, ZN => n6376);
   U4136 : NAND2_X1 port map( A1 => n6377, A2 => n6376, ZN => n6379);
   U4137 : INV_X1 port map( A => n6379, ZN => n6378);
   U4138 : NAND2_X1 port map( A1 => n6380, A2 => n6379, ZN => n6406);
   U4140 : INV_X1 port map( A => n6382, ZN => n6383);
   U4141 : AOI21_X1 port map( B1 => n8549, B2 => n6383, A => n4975, ZN => n6405
                           );
   U4142 : MUX2_X1 port map( A => n7123, B => n7122, S => n377, Z => n6387);
   U4143 : XNOR2_X1 port map( A => n8403, B => n360, ZN => n6385);
   U4144 : NAND2_X1 port map( A1 => n5307, A2 => n6385, ZN => n6386);
   U4145 : NAND2_X1 port map( A1 => n6387, A2 => n6386, ZN => n6413);
   U4146 : INV_X1 port map( A => n6409, ZN => n6414);
   U4147 : XNOR2_X1 port map( A => n6413, B => n6414, ZN => n6390);
   U4148 : MUX2_X1 port map( A => n8445, B => n6740, S => n357, Z => n6412);
   U4149 : MUX2_X1 port map( A => n8459, B => n8434, S => n8334, Z => n6411);
   U4150 : NAND2_X1 port map( A1 => n6412, A2 => n6411, ZN => n6389);
   U4151 : XNOR2_X1 port map( A => n6390, B => n6389, ZN => n6421);
   U4152 : OAI21_X1 port map( B1 => n6391, B2 => n6419, A => n6421, ZN => n6393
                           );
   U4153 : NAND2_X1 port map( A1 => n6391, A2 => n6419, ZN => n6392);
   U4154 : NAND2_X1 port map( A1 => n6393, A2 => n6392, ZN => n6661);
   U4155 : INV_X1 port map( A => n6395, ZN => n6404);
   U4156 : NAND2_X1 port map( A1 => n6395, A2 => n6394, ZN => n6402);
   U4157 : AND3_X1 port map( A1 => n6398, A2 => n6397, A3 => n6396, ZN => n6400
                           );
   U4158 : NAND2_X1 port map( A1 => n6400, A2 => n6399, ZN => n6401);
   U4159 : NAND2_X1 port map( A1 => n6406, A2 => n6405, ZN => n6408);
   U4160 : NAND2_X1 port map( A1 => n6408, A2 => n6407, ZN => n6645);
   U4163 : INV_X1 port map( A => n6413, ZN => n6415);
   U4164 : NAND2_X1 port map( A1 => n6415, A2 => n6414, ZN => n6416);
   U4165 : NAND2_X1 port map( A1 => n6417, A2 => n6416, ZN => n6646);
   U4166 : XNOR2_X1 port map( A => n6661, B => n6660, ZN => n6418);
   U4167 : XNOR2_X1 port map( A => n6664, B => n6418, ZN => n6669);
   U4168 : XNOR2_X1 port map( A => n6668, B => n6669, ZN => n6488);
   U4169 : XNOR2_X1 port map( A => n6420, B => n4403, ZN => n6423);
   U4170 : INV_X1 port map( A => n6421, ZN => n6422);
   U4171 : XNOR2_X1 port map( A => n6423, B => n6422, ZN => n6578);
   U4172 : INV_X1 port map( A => n6424, ZN => n6429);
   U4173 : INV_X1 port map( A => n6427, ZN => n6425);
   U4174 : INV_X1 port map( A => n8429, ZN => n6428);
   U4175 : NAND2_X1 port map( A1 => n6430, A2 => n4892, ZN => n6433);
   U4177 : AOI22_X1 port map( A1 => n6434, A2 => n6433, B1 => n8415, B2 => 
                           n6431, ZN => n6435);
   U4178 : NAND2_X1 port map( A1 => n6436, A2 => n8565, ZN => n6482);
   U4179 : NAND2_X1 port map( A1 => n6482, A2 => n6483, ZN => n6441);
   U4180 : INV_X1 port map( A => n6437, ZN => n6439);
   U4181 : OAI21_X1 port map( B1 => n6440, B2 => n6439, A => n6438, ZN => n6653
                           );
   U4182 : NAND2_X1 port map( A1 => n6578, A2 => n8566, ZN => n6569);
   U4183 : INV_X1 port map( A => n6442, ZN => n6446);
   U4185 : OAI21_X1 port map( B1 => n6446, B2 => n6445, A => n8548, ZN => n6448
                           );
   U4186 : NAND2_X1 port map( A1 => n6446, A2 => n6445, ZN => n6447);
   U4187 : NAND2_X1 port map( A1 => n6448, A2 => n6447, ZN => n6573);
   U4188 : NAND2_X1 port map( A1 => n6569, A2 => n6573, ZN => n6450);
   U4189 : INV_X1 port map( A => n6578, ZN => n6449);
   U4190 : INV_X1 port map( A => n6493, ZN => n6574);
   U4191 : NAND2_X1 port map( A1 => n6449, A2 => n6574, ZN => n6568);
   U4192 : NAND2_X1 port map( A1 => n6450, A2 => n6568, ZN => n6487);
   U4193 : INV_X1 port map( A => n6451, ZN => n6453);
   U4194 : OAI21_X1 port map( B1 => n6454, B2 => n6453, A => n6452, ZN => n6456
                           );
   U4195 : NAND2_X1 port map( A1 => n6454, A2 => n6453, ZN => n6455);
   U4196 : NAND2_X1 port map( A1 => n6456, A2 => n6455, ZN => n6570);
   U4197 : XNOR2_X1 port map( A => A_SIG_23_port, B => n362, ZN => n6457);
   U4198 : NAND2_X1 port map( A1 => n6457, A2 => n5749, ZN => n6458);
   U4199 : INV_X1 port map( A => n6469, ZN => n6466);
   U4200 : NAND2_X1 port map( A1 => n6460, A2 => n8394, ZN => n6462);
   U4201 : NAND2_X1 port map( A1 => n5226, A2 => n359, ZN => n6461);
   U4202 : NAND2_X1 port map( A1 => n6462, A2 => n6461, ZN => n6465);
   U4203 : XNOR2_X1 port map( A => n377, B => n6229, ZN => n6463);
   U4204 : NOR2_X1 port map( A1 => n6687, A2 => n6463, ZN => n6464);
   U4205 : NOR2_X1 port map( A1 => n6465, A2 => n6464, ZN => n6467);
   U4206 : NAND2_X1 port map( A1 => n6466, A2 => n6467, ZN => n6584);
   U4208 : NAND2_X1 port map( A1 => n6469, A2 => n8481, ZN => n6583);
   U4209 : NAND2_X1 port map( A1 => n6584, A2 => n6583, ZN => n6472);
   U4210 : MUX2_X1 port map( A => n6714, B => n6888, S => n205, Z => n6471);
   U4211 : MUX2_X1 port map( A => n6715, B => n6887, S => n8423, Z => n6470);
   U4212 : NAND2_X1 port map( A1 => n6471, A2 => n6470, ZN => n6585);
   U4213 : XNOR2_X1 port map( A => n6472, B => n6585, ZN => n6650);
   U4214 : NAND2_X1 port map( A1 => n6476, A2 => n6477, ZN => n6473);
   U4215 : NAND3_X1 port map( A1 => n6475, A2 => n6474, A3 => n6473, ZN => 
                           n6481);
   U4216 : INV_X1 port map( A => n6476, ZN => n6479);
   U4217 : INV_X1 port map( A => n6477, ZN => n6478);
   U4218 : NAND2_X1 port map( A1 => n6479, A2 => n6478, ZN => n6480);
   U4219 : NAND2_X1 port map( A1 => n6481, A2 => n6480, ZN => n6656);
   U4220 : XNOR2_X1 port map( A => n6650, B => n6656, ZN => n6485);
   U4221 : NAND2_X1 port map( A1 => n6482, A2 => n6653, ZN => n6484);
   U4222 : NAND2_X1 port map( A1 => n6484, A2 => n6483, ZN => n6652);
   U4223 : XNOR2_X1 port map( A => n6485, B => n6652, ZN => n6572);
   U4224 : XNOR2_X1 port map( A => n6572, B => n6570, ZN => n6486);
   U4225 : XNOR2_X1 port map( A => n6487, B => n6486, ZN => n6670);
   U4227 : NAND2_X1 port map( A1 => n6489, A2 => n6490, ZN => n6492);
   U4228 : INV_X1 port map( A => n6548, ZN => n6491);
   U4229 : XNOR2_X1 port map( A => n6492, B => n6491, ZN => n6513);
   U4230 : XNOR2_X1 port map( A => n6493, B => n6573, ZN => n6494);
   U4231 : XNOR2_X1 port map( A => n6578, B => n6494, ZN => n6546);
   U4232 : XNOR2_X1 port map( A => n6496, B => n6495, ZN => n6498);
   U4233 : XNOR2_X1 port map( A => n6498, B => n6497, ZN => n6529);
   U4235 : AOI21_X1 port map( B1 => n6500, B2 => n6501, A => n6499, ZN => n6528
                           );
   U4236 : NAND2_X1 port map( A1 => n6506, A2 => n6503, ZN => n6505);
   U4237 : NAND2_X1 port map( A1 => n6504, A2 => n6505, ZN => n6510);
   U4239 : NAND2_X1 port map( A1 => n8573, A2 => n6507, ZN => n6509);
   U4240 : NAND2_X1 port map( A1 => n6510, A2 => n6509, ZN => n6531);
   U4241 : FA_X1 port map( A => n8574, B => n6502, CI => n6531, CO => n6552, S 
                           => n_1140);
   U4242 : OAI21_X1 port map( B1 => n6513, B2 => n6512, A => n6552, ZN => n6515
                           );
   U4243 : NAND2_X1 port map( A1 => n6513, A2 => n6512, ZN => n6514);
   U4244 : NAND2_X1 port map( A1 => n6515, A2 => n6514, ZN => n6561);
   U4246 : NAND2_X1 port map( A1 => n8073, A2 => n8484, ZN => n7651);
   U4247 : NAND2_X1 port map( A1 => n6517, A2 => n6516, ZN => n6540);
   U4248 : NAND2_X1 port map( A1 => n6541, A2 => n6540, ZN => n6518);
   U4249 : XNOR2_X1 port map( A => n6518, B => n6539, ZN => n6519);
   U4250 : NAND2_X1 port map( A1 => n6519, A2 => n6524, ZN => n6527);
   U4252 : OAI21_X1 port map( B1 => n6525, B2 => n6524, A => n6523, ZN => n6526
                           );
   U4253 : NAND2_X1 port map( A1 => n6527, A2 => n6526, ZN => n6563);
   U4254 : INV_X1 port map( A => n6528, ZN => n6530);
   U4255 : XNOR2_X1 port map( A => n6530, B => n6529, ZN => n6533);
   U4256 : INV_X1 port map( A => n6531, ZN => n6532);
   U4258 : INV_X1 port map( A => n6534, ZN => n6535);
   U4259 : XNOR2_X1 port map( A => n6536, B => n6535, ZN => n6537);
   U4260 : XNOR2_X1 port map( A => n6538, B => n6537, ZN => n6556);
   U4261 : XNOR2_X1 port map( A => n4413, B => n6556, ZN => n6543);
   U4262 : NAND2_X1 port map( A1 => n6540, A2 => n6539, ZN => n6542);
   U4263 : NAND2_X1 port map( A1 => n6542, A2 => n6541, ZN => n6558);
   U4264 : XNOR2_X1 port map( A => n6543, B => n8534, ZN => n6564);
   U4265 : NAND2_X1 port map( A1 => n4492, A2 => n4431, ZN => n8057);
   U4266 : INV_X1 port map( A => n6544, ZN => n6545);
   U4267 : XNOR2_X1 port map( A => n6546, B => n6545, ZN => n6551);
   U4268 : INV_X1 port map( A => n6547, ZN => n6549);
   U4269 : XNOR2_X1 port map( A => n6549, B => n6548, ZN => n6550);
   U4270 : XNOR2_X1 port map( A => n6551, B => n6550, ZN => n6554);
   U4271 : INV_X1 port map( A => n6552, ZN => n6553);
   U4272 : NAND2_X1 port map( A1 => n8077, A2 => n4444, ZN => n8074);
   U4273 : NAND2_X1 port map( A1 => n8057, A2 => n8558, ZN => n7650);
   U4275 : INV_X1 port map( A => n8096, ZN => n6566);
   U4276 : INV_X1 port map( A => n7623, ZN => n6560);
   U4277 : NAND2_X1 port map( A1 => n6560, A2 => n8484, ZN => n7735);
   U4278 : INV_X1 port map( A => n8086, ZN => n6562);
   U4279 : INV_X1 port map( A => n6561, ZN => n8085);
   U4280 : NAND2_X1 port map( A1 => n6562, A2 => n8085, ZN => n7734);
   U4281 : AND2_X1 port map( A1 => n7735, A2 => n7734, ZN => n7595);
   U4282 : AND2_X1 port map( A1 => n6564, A2 => n6563, ZN => n8079);
   U4283 : NAND3_X1 port map( A1 => n8079, A2 => n8586, A3 => n8542, ZN => 
                           n6565);
   U4284 : NAND2_X1 port map( A1 => n7595, A2 => n6565, ZN => n8100);
   U4285 : AOI21_X1 port map( B1 => n8444, B2 => n6566, A => n8100, ZN => n6676
                           );
   U4286 : INV_X1 port map( A => n6573, ZN => n6567);
   U4287 : NAND2_X1 port map( A1 => n6568, A2 => n6567, ZN => n6582);
   U4288 : INV_X1 port map( A => n6570, ZN => n6581);
   U4289 : NAND2_X1 port map( A1 => n6572, A2 => n6569, ZN => n6571);
   U4290 : NAND2_X1 port map( A1 => n6571, A2 => n6570, ZN => n6580);
   U4291 : NOR2_X1 port map( A1 => n6574, A2 => n6573, ZN => n6577);
   U4292 : INV_X1 port map( A => n6572, ZN => n6576);
   U4293 : NAND2_X1 port map( A1 => n6574, A2 => n6573, ZN => n6575);
   U4294 : OAI211_X1 port map( C1 => n6578, C2 => n6577, A => n6576, B => n6575
                           , ZN => n6579);
   U4295 : OAI211_X1 port map( C1 => n6582, C2 => n6581, A => n6580, B => n6579
                           , ZN => n6776);
   U4296 : INV_X1 port map( A => n6583, ZN => n6586);
   U4297 : MUX2_X1 port map( A => n6800, B => n7508, S => n379, Z => n6597);
   U4298 : XNOR2_X1 port map( A => n4381, B => n6593, ZN => n6594);
   U4299 : NAND2_X1 port map( A1 => n6594, A2 => n6595, ZN => n6596);
   U4300 : NAND2_X1 port map( A1 => n6597, A2 => n6596, ZN => n6742);
   U4301 : NAND2_X1 port map( A1 => A_SIG_23_port, A2 => n8352, ZN => n6846);
   U4302 : XNOR2_X1 port map( A => n8560, B => n6846, ZN => n6600);
   U4303 : NAND2_X1 port map( A1 => n6740, A2 => n8434, ZN => n6598);
   U4304 : AOI21_X1 port map( B1 => n8397, B2 => n8335, A => n8002, ZN => n6843
                           );
   U4305 : MUX2_X1 port map( A => n6598, B => n6843, S => n7506, Z => n6599);
   U4306 : XNOR2_X1 port map( A => n6600, B => n6599, ZN => n6931);
   U4307 : INV_X1 port map( A => n6602, ZN => n6950);
   U4308 : INV_X1 port map( A => n6948, ZN => n6951);
   U4311 : INV_X1 port map( A => n6605, ZN => n6612);
   U4312 : NAND2_X1 port map( A1 => n8324, A2 => n376, ZN => n6609);
   U4313 : MUX2_X1 port map( A => n7692, B => n7254, S => n8333, Z => n6613);
   U4314 : INV_X1 port map( A => n7690, ZN => n7392);
   U4315 : NAND2_X1 port map( A1 => n6617, A2 => n6616, ZN => n6723);
   U4316 : NAND2_X1 port map( A1 => n6723, A2 => n6721, ZN => n6623);
   U4317 : NAND3_X1 port map( A1 => n6620, A2 => n6619, A3 => n6618, ZN => 
                           n6622);
   U4318 : NAND2_X1 port map( A1 => n6622, A2 => n6621, ZN => n6722);
   U4319 : XNOR2_X1 port map( A => n6624, B => n6958, ZN => n6625);
   U4320 : XNOR2_X1 port map( A => n6682, B => n6625, ZN => n6777);
   U4321 : XNOR2_X1 port map( A => n6776, B => n6777, ZN => n6667);
   U4322 : MUX2_X1 port map( A => n7195, B => n7080, S => n360, Z => n6627);
   U4323 : MUX2_X1 port map( A => n7324, B => n7323, S => n8332, Z => n6626);
   U4324 : NAND2_X1 port map( A1 => n6627, A2 => n6626, ZN => n6753);
   U4325 : MUX2_X1 port map( A => n4490, B => n7084, S => n8423, Z => n6629);
   U4326 : MUX2_X1 port map( A => n4607, B => n8596, S => n371, Z => n6628);
   U4327 : NAND2_X1 port map( A1 => n6629, A2 => n6628, ZN => n6754);
   U4328 : XNOR2_X1 port map( A => n6754, B => n6753, ZN => n6632);
   U4329 : MUX2_X1 port map( A => n8501, B => n7053, S => n359, Z => n6631);
   U4330 : MUX2_X1 port map( A => n4462, B => n7054, S => n8326, Z => n6630);
   U4331 : NAND2_X1 port map( A1 => n6631, A2 => n6630, ZN => n6757);
   U4332 : XNOR2_X1 port map( A => n6632, B => n6757, ZN => n6640);
   U4333 : MUX2_X1 port map( A => n7086, B => n7047, S => n204, Z => n6634);
   U4334 : MUX2_X1 port map( A => n8559, B => n8582, S => n8327, Z => n6633);
   U4335 : NAND2_X1 port map( A1 => n6634, A2 => n6633, ZN => n6764);
   U4336 : MUX2_X1 port map( A => n6811, B => n4360, S => n363, Z => n6636);
   U4337 : MUX2_X1 port map( A => n7123, B => n6812, S => n372, Z => n6635);
   U4338 : NAND2_X1 port map( A1 => n6636, A2 => n6635, ZN => n6763);
   U4339 : XNOR2_X1 port map( A => n6763, B => n6764, ZN => n6639);
   U4340 : MUX2_X1 port map( A => n6714, B => n6888, S => n357, Z => n6638);
   U4341 : MUX2_X1 port map( A => n6715, B => n6243, S => n205, Z => n6637);
   U4342 : NAND2_X1 port map( A1 => n6638, A2 => n6637, ZN => n6760);
   U4343 : XNOR2_X1 port map( A => n6639, B => n6760, ZN => n6641);
   U4344 : NAND2_X1 port map( A1 => n6640, A2 => n6641, ZN => n6728);
   U4345 : INV_X1 port map( A => n6640, ZN => n6643);
   U4346 : INV_X1 port map( A => n6641, ZN => n6642);
   U4347 : NAND2_X1 port map( A1 => n6643, A2 => n6642, ZN => n6729);
   U4348 : NAND2_X1 port map( A1 => n6728, A2 => n6729, ZN => n6649);
   U4349 : OAI21_X1 port map( B1 => n6647, B2 => n6646, A => n6645, ZN => n6731
                           );
   U4350 : NAND2_X1 port map( A1 => n6647, A2 => n6646, ZN => n6726);
   U4351 : NAND2_X1 port map( A1 => n6731, A2 => n6726, ZN => n6648);
   U4352 : XNOR2_X1 port map( A => n6649, B => n6648, ZN => n6681);
   U4353 : INV_X1 port map( A => n6650, ZN => n6651);
   U4354 : OAI21_X1 port map( B1 => n6652, B2 => n6656, A => n6651, ZN => n6658
                           );
   U4355 : INV_X1 port map( A => n6653, ZN => n6654);
   U4356 : NAND2_X1 port map( A1 => n6483, A2 => n6654, ZN => n6655);
   U4357 : NAND3_X1 port map( A1 => n6656, A2 => n6655, A3 => n6482, ZN => 
                           n6657);
   U4358 : NAND2_X1 port map( A1 => n6658, A2 => n6657, ZN => n6677);
   U4359 : XNOR2_X1 port map( A => n6681, B => n6677, ZN => n6666);
   U4360 : INV_X1 port map( A => n6661, ZN => n6665);
   U4361 : INV_X1 port map( A => n6660, ZN => n6659);
   U4362 : OR2_X1 port map( A1 => n6664, A2 => n6659, ZN => n6663);
   U4363 : NAND2_X1 port map( A1 => n6661, A2 => n6660, ZN => n6662);
   U4364 : XNOR2_X1 port map( A => n4429, B => n6666, ZN => n6778);
   U4365 : XNOR2_X1 port map( A => n6667, B => n6778, ZN => n7492);
   U4366 : INV_X1 port map( A => n6669, ZN => n6671);
   U4367 : OAI21_X1 port map( B1 => n4476, B2 => n6671, A => n6670, ZN => n6673
                           );
   U4368 : NAND2_X1 port map( A1 => n4476, A2 => n6671, ZN => n6672);
   U4369 : NAND2_X1 port map( A1 => n6673, A2 => n6672, ZN => n8098);
   U4370 : XNOR2_X1 port map( A => n8584, B => n8098, ZN => n6675);
   U4371 : NAND2_X1 port map( A1 => n6676, A2 => n6675, ZN => n6674);
   U4372 : OAI21_X1 port map( B1 => n6675, B2 => n6676, A => n6674, ZN => 
                           I2_dtemp_30_port);
   U4373 : INV_X1 port map( A => n8536, ZN => n6679);
   U4374 : INV_X1 port map( A => n6677, ZN => n6678);
   U4375 : AOI21_X1 port map( B1 => n6680, B2 => n6679, A => n6678, ZN => n6979
                           );
   U4376 : AND2_X1 port map( A1 => n4429, A2 => n8536, ZN => n6980);
   U4377 : OAI21_X1 port map( B1 => n4421, B2 => n6958, A => n6959, ZN => n6684
                           );
   U4378 : NAND2_X1 port map( A1 => n4421, A2 => n6958, ZN => n6683);
   U4379 : NAND2_X1 port map( A1 => n6684, A2 => n6683, ZN => n6947);
   U4380 : XNOR2_X1 port map( A => n372, B => n6229, ZN => n6686);
   U4381 : NOR2_X1 port map( A1 => n6687, A2 => n6686, ZN => n6692);
   U4382 : NAND2_X1 port map( A1 => n5226, A2 => n360, ZN => n6689);
   U4383 : NAND2_X1 port map( A1 => n6689, A2 => n6690, ZN => n6691);
   U4384 : INV_X1 port map( A => n6843, ZN => n6838);
   U4385 : XNOR2_X1 port map( A => n6839, B => n6838, ZN => n6695);
   U4386 : MUX2_X1 port map( A => n6811, B => n4360, S => n371, Z => n6694);
   U4388 : NAND2_X1 port map( A1 => n6694, A2 => n6693, ZN => n6842);
   U4389 : XNOR2_X1 port map( A => n6842, B => n6695, ZN => n6719);
   U4390 : MUX2_X1 port map( A => n7090, B => n8581, S => n204, Z => n6700);
   U4391 : XNOR2_X1 port map( A => n8503, B => n8392, ZN => n6698);
   U4392 : NAND2_X1 port map( A1 => n6374, A2 => n6698, ZN => n6699);
   U4393 : NAND2_X1 port map( A1 => n6700, A2 => n6699, ZN => n6713);
   U4394 : XNOR2_X1 port map( A => n8353, B => n377, ZN => n6701);
   U4395 : NAND2_X1 port map( A1 => n6702, A2 => n6701, ZN => n6711);
   U4398 : NAND3_X1 port map( A1 => n8369, A2 => n8394, A3 => n6705, ZN => 
                           n6707);
   U4399 : NAND2_X1 port map( A1 => n6707, A2 => n6706, ZN => n6708);
   U4400 : NAND2_X1 port map( A1 => n6709, A2 => n6708, ZN => n6710);
   U4401 : NAND2_X1 port map( A1 => n6711, A2 => n6710, ZN => n6712);
   U4402 : NAND2_X1 port map( A1 => n6713, A2 => n6712, ZN => n6855);
   U4403 : NAND2_X1 port map( A1 => n6853, A2 => n6855, ZN => n6718);
   U4404 : MUX2_X1 port map( A => n6714, B => n6888, S => n7506, Z => n6717);
   U4405 : MUX2_X1 port map( A => n6715, B => n6243, S => n357, Z => n6716);
   U4406 : XNOR2_X1 port map( A => n6718, B => n6852, ZN => n6720);
   U4407 : NAND2_X1 port map( A1 => n6720, A2 => n6719, ZN => n6919);
   U4408 : NAND2_X1 port map( A1 => n6921, A2 => n6919, ZN => n6725);
   U4409 : NAND2_X1 port map( A1 => n6721, A2 => n6722, ZN => n6724);
   U4410 : NAND2_X1 port map( A1 => n6724, A2 => n6723, ZN => n6920);
   U4411 : XNOR2_X1 port map( A => n6725, B => n6920, ZN => n6946);
   U4412 : INV_X1 port map( A => n6946, ZN => n6957);
   U4413 : INV_X1 port map( A => n6728, ZN => n6732);
   U4414 : INV_X1 port map( A => n6726, ZN => n6727);
   U4415 : NAND2_X1 port map( A1 => n4425, A2 => n6727, ZN => n6730);
   U4416 : OAI211_X1 port map( C1 => n6732, C2 => n6731, A => n6729, B => n6730
                           , ZN => n6962);
   U4417 : XNOR2_X1 port map( A => n6962, B => n6957, ZN => n6733);
   U4418 : XNOR2_X1 port map( A => n6733, B => n6947, ZN => n6775);
   U4419 : INV_X1 port map( A => n8599, ZN => n6737);
   U4420 : INV_X1 port map( A => n8587, ZN => n6736);
   U4421 : AOI21_X1 port map( B1 => n6737, B2 => n6931, A => n6736, ZN => n6911
                           );
   U4422 : AND2_X1 port map( A1 => n8599, A2 => n4406, ZN => n6910);
   U4424 : AOI21_X1 port map( B1 => n6738, B2 => n7506, A => n6846, ZN => n6739
                           );
   U4425 : OAI211_X1 port map( C1 => n7769, C2 => n8434, A => n6740, B => n6739
                           , ZN => n6741);
   U4426 : NAND2_X1 port map( A1 => n6742, A2 => n6741, ZN => n6747);
   U4427 : AOI22_X1 port map( A1 => n8434, A2 => n8336, B1 => n7506, B2 => 
                           n6743, ZN => n6745);
   U4428 : OAI21_X1 port map( B1 => n6745, B2 => n6744, A => n6846, ZN => n6746
                           );
   U4429 : NAND2_X1 port map( A1 => n6747, A2 => n6746, ZN => n6860);
   U4430 : MUX2_X1 port map( A => n7253, B => n7392, S => n8327, Z => n6749);
   U4431 : MUX2_X1 port map( A => n7692, B => n7773, S => n7945, Z => n6748);
   U4432 : NAND2_X1 port map( A1 => n6749, A2 => n6748, ZN => n6859);
   U4433 : XNOR2_X1 port map( A => n6860, B => n6859, ZN => n6752);
   U4434 : MUX2_X1 port map( A => n4490, B => n7051, S => n205, Z => n6751);
   U4435 : MUX2_X1 port map( A => n4607, B => n8596, S => n8423, Z => n6750);
   U4436 : NAND2_X1 port map( A1 => n6751, A2 => n6750, ZN => n6858);
   U4438 : XNOR2_X1 port map( A => n8576, B => n6935, ZN => n6773);
   U4439 : NAND2_X1 port map( A1 => n6753, A2 => n6757, ZN => n6756);
   U4441 : NAND2_X1 port map( A1 => n6756, A2 => n8448, ZN => n6759);
   U4442 : NAND2_X1 port map( A1 => n6759, A2 => n6758, ZN => n6864);
   U4443 : INV_X1 port map( A => n6864, ZN => n6772);
   U4444 : INV_X1 port map( A => n6760, ZN => n6762);
   U4445 : NAND2_X1 port map( A1 => n6764, A2 => n6763, ZN => n6761);
   U4446 : NAND2_X1 port map( A1 => n6762, A2 => n6761, ZN => n6767);
   U4447 : INV_X1 port map( A => n6764, ZN => n6765);
   U4448 : NAND2_X1 port map( A1 => n4436, A2 => n6765, ZN => n6766);
   U4449 : NAND2_X1 port map( A1 => n6767, A2 => n6766, ZN => n6862);
   U4450 : MUX2_X1 port map( A => n8476, B => n7559, S => n356, Z => n6769);
   U4451 : MUX2_X1 port map( A => n7227, B => n7439, S => n373, Z => n6768);
   U4452 : NAND2_X1 port map( A1 => n6769, A2 => n6768, ZN => n6851);
   U4453 : INV_X1 port map( A => n6846, ZN => n6849);
   U4454 : NAND2_X1 port map( A1 => A_SIG_23_port, A2 => n8333, ZN => n6847);
   U4455 : XNOR2_X1 port map( A => n6849, B => n6847, ZN => n6770);
   U4456 : XNOR2_X1 port map( A => n6851, B => n6770, ZN => n6863);
   U4457 : XNOR2_X1 port map( A => n6862, B => n6863, ZN => n6771);
   U4458 : XNOR2_X1 port map( A => n8589, B => n6772, ZN => n6915);
   U4459 : XNOR2_X1 port map( A => n6773, B => n4456, ZN => n6774);
   U4460 : NAND2_X1 port map( A1 => n6775, A2 => n6774, ZN => n6981);
   U4461 : NAND2_X1 port map( A1 => n6778, A2 => n6777, ZN => n6779);
   U4462 : INV_X1 port map( A => n8123, ZN => n8111);
   U4463 : NAND2_X1 port map( A1 => n7253, A2 => n8351, ZN => n6781);
   U4464 : OAI21_X1 port map( B1 => n7690, B2 => n8351, A => n6781, ZN => n6783
                           );
   U4465 : MUX2_X1 port map( A => n7692, B => n7254, S => B_SIG_9_port, Z => 
                           n6782);
   U4466 : MUX2_X1 port map( A => n7195, B => n7080, S => n363, Z => n6785);
   U4467 : MUX2_X1 port map( A => n7324, B => n7323, S => n8330, Z => n6784);
   U4468 : NAND2_X1 port map( A1 => n6785, A2 => n6784, ZN => n7023);
   U4469 : NAND2_X1 port map( A1 => n7021, A2 => n7023, ZN => n6788);
   U4470 : MUX2_X1 port map( A => n8501, B => n7053, S => n360, Z => n6787);
   U4471 : MUX2_X1 port map( A => n4461, B => n7054, S => n8332, Z => n6786);
   U4473 : NAND2_X1 port map( A1 => n6788, A2 => n7022, ZN => n6792);
   U4475 : INV_X1 port map( A => n4486, ZN => n6789);
   U4476 : NAND2_X1 port map( A1 => n8472, A2 => n6789, ZN => n6791);
   U4477 : NAND2_X1 port map( A1 => n6792, A2 => n6791, ZN => n6797);
   U4478 : MUX2_X1 port map( A => n6811, B => n7120, S => n205, Z => n6794);
   U4479 : MUX2_X1 port map( A => n7123, B => n7122, S => n8423, Z => n6793);
   U4480 : NAND2_X1 port map( A1 => n6793, A2 => n6794, ZN => n7043);
   U4481 : AND2_X1 port map( A1 => B_SIG_8_port, A2 => A_SIG_23_port, ZN => 
                           n6808);
   U4482 : INV_X1 port map( A => n6808, ZN => n6809);
   U4483 : NAND2_X1 port map( A1 => B_SIG_9_port, A2 => n8504, ZN => n6795);
   U4484 : OR2_X1 port map( A1 => n6809, A2 => n6795, ZN => n7044);
   U4485 : NAND2_X1 port map( A1 => n6809, A2 => n6795, ZN => n7042);
   U4486 : NAND2_X1 port map( A1 => n7044, A2 => n7042, ZN => n6796);
   U4487 : XNOR2_X1 port map( A => n7043, B => n6796, ZN => n7020);
   U4488 : XNOR2_X1 port map( A => n6797, B => n7020, ZN => n6806);
   U4489 : MUX2_X1 port map( A => n7195, B => n7080, S => n371, Z => n6799);
   U4490 : MUX2_X1 port map( A => n7324, B => n8465, S => n8329, Z => n6798);
   U4491 : NAND2_X1 port map( A1 => n6799, A2 => n6798, ZN => n6998);
   U4492 : MUX2_X1 port map( A => n5866, B => n5867, S => n377, Z => n6802);
   U4493 : MUX2_X1 port map( A => n6800, B => n7508, S => n359, Z => n6801);
   U4494 : NAND2_X1 port map( A1 => n6802, A2 => n6801, ZN => n6996);
   U4495 : XNOR2_X1 port map( A => n6996, B => n6998, ZN => n6805);
   U4496 : MUX2_X1 port map( A => n8500, B => n7053, S => n372, Z => n6804);
   U4497 : MUX2_X1 port map( A => n4462, B => n7054, S => n8337, Z => n6803);
   U4498 : XNOR2_X1 port map( A => n6805, B => n7001, ZN => n7027);
   U4499 : XNOR2_X1 port map( A => n7027, B => n6806, ZN => n6837);
   U4501 : MUX2_X1 port map( A => n7094, B => n7093, S => n359, Z => n6807);
   U4502 : NAND2_X1 port map( A1 => n6810, A2 => n6808, ZN => n6883);
   U4503 : OR2_X1 port map( A1 => n6810, A2 => n6808, ZN => n6881);
   U4504 : NAND2_X1 port map( A1 => n6883, A2 => n6881, ZN => n6816);
   U4505 : MUX2_X1 port map( A => n7123, B => n7122, S => n371, Z => n6814);
   U4506 : NAND2_X1 port map( A1 => n6815, A2 => n6814, ZN => n6882);
   U4507 : XNOR2_X1 port map( A => n6816, B => n6882, ZN => n6916);
   U4508 : INV_X1 port map( A => n6817, ZN => n6818);
   U4509 : MUX2_X1 port map( A => n6819, B => n6818, S => n7769, Z => n6820);
   U4510 : NAND2_X1 port map( A1 => n6820, A2 => n6888, ZN => n6875);
   U4511 : NAND2_X1 port map( A1 => n8469, A2 => n8334, ZN => n6822);
   U4512 : NAND2_X1 port map( A1 => n6822, A2 => n6821, ZN => n6825);
   U4513 : XNOR2_X1 port map( A => n8331, B => n5883, ZN => n6823);
   U4514 : NAND2_X1 port map( A1 => n4491, A2 => n6823, ZN => n6824);
   U4515 : NAND2_X1 port map( A1 => n6825, A2 => n6824, ZN => n6874);
   U4516 : XNOR2_X1 port map( A => n6874, B => n6875, ZN => n6828);
   U4517 : MUX2_X1 port map( A => n7047, B => n7086, S => n4381, Z => n6827);
   U4518 : MUX2_X1 port map( A => n8559, B => n8582, S => n379, Z => n6826);
   U4519 : NAND2_X1 port map( A1 => n6827, A2 => n6826, ZN => n6876);
   U4520 : XNOR2_X1 port map( A => n6876, B => n6828, ZN => n6917);
   U4521 : NAND2_X1 port map( A1 => n6916, A2 => n6917, ZN => n6830);
   U4522 : XNOR2_X1 port map( A => n7023, B => n7021, ZN => n6829);
   U4523 : XNOR2_X1 port map( A => n6829, B => n7022, ZN => n6918);
   U4524 : NAND2_X1 port map( A1 => n6830, A2 => n6918, ZN => n6834);
   U4525 : INV_X1 port map( A => n8554, ZN => n6832);
   U4526 : INV_X1 port map( A => n6917, ZN => n6831);
   U4527 : NAND2_X1 port map( A1 => n6832, A2 => n6831, ZN => n6833);
   U4528 : NAND2_X1 port map( A1 => n6834, A2 => n6833, ZN => n6836);
   U4529 : NAND2_X1 port map( A1 => n8551, A2 => n6836, ZN => n6992);
   U4531 : AND2_X1 port map( A1 => n6994, A2 => n6992, ZN => n6873);
   U4532 : NAND2_X1 port map( A1 => n4473, A2 => n6838, ZN => n6841);
   U4534 : NAND2_X1 port map( A1 => n8474, A2 => n6844, ZN => n6868);
   U4535 : NOR2_X1 port map( A1 => n6846, A2 => n6847, ZN => n6850);
   U4536 : INV_X1 port map( A => n6847, ZN => n6848);
   U4537 : XNOR2_X1 port map( A => n6868, B => n6867, ZN => n6857);
   U4538 : XNOR2_X1 port map( A => n6857, B => n6869, ZN => n6861);
   U4539 : FA_X1 port map( A => n6859, B => n6860, CI => n6858, CO => n6870, S 
                           => n_1141);
   U4540 : NAND2_X1 port map( A1 => n6861, A2 => n6870, ZN => n6941);
   U4541 : OAI21_X1 port map( B1 => n6864, B2 => n8588, A => n6862, ZN => n6866
                           );
   U4542 : NAND2_X1 port map( A1 => n6864, A2 => n8588, ZN => n6865);
   U4543 : NAND2_X1 port map( A1 => n6866, A2 => n6865, ZN => n6943);
   U4544 : NAND2_X1 port map( A1 => n6941, A2 => n6943, ZN => n6872);
   U4545 : NAND2_X1 port map( A1 => n4440, A2 => n6867, ZN => n6903);
   U4546 : INV_X1 port map( A => n6869, ZN => n6906);
   U4547 : INV_X1 port map( A => n6870, ZN => n6871);
   U4548 : NAND2_X1 port map( A1 => n6872, A2 => n6942, ZN => n6995);
   U4549 : XNOR2_X1 port map( A => n6873, B => n6995, ZN => n6909);
   U4550 : AOI21_X1 port map( B1 => n6876, B2 => n6875, A => n6874, ZN => n6878
                           );
   U4551 : NOR2_X1 port map( A1 => n6876, A2 => n6875, ZN => n6877);
   U4552 : MUX2_X1 port map( A => n7253, B => n7771, S => n379, Z => n6880);
   U4553 : MUX2_X1 port map( A => n7692, B => n7773, S => n8351, Z => n6879);
   U4554 : NAND2_X1 port map( A1 => n6880, A2 => n6879, ZN => n6896);
   U4555 : NAND2_X1 port map( A1 => n6895, A2 => n6896, ZN => n7061);
   U4556 : NAND2_X1 port map( A1 => n7061, A2 => n7060, ZN => n6884);
   U4557 : XNOR2_X1 port map( A => n6884, B => n6898, ZN => n6894);
   U4558 : MUX2_X1 port map( A => n7665, B => n7556, S => n356, Z => n6886);
   U4559 : MUX2_X1 port map( A => n7696, B => n7695, S => n373, Z => n6885);
   U4560 : NAND2_X1 port map( A1 => n6886, A2 => n6885, ZN => n7005);
   U4561 : AND2_X1 port map( A1 => n6888, A2 => n6887, ZN => n7006);
   U4562 : XNOR2_X1 port map( A => n7005, B => n7006, ZN => n6893);
   U4563 : MUX2_X1 port map( A => n4489, B => n7084, S => n7506, Z => n6892);
   U4564 : MUX2_X1 port map( A => n8469, B => n8595, S => n357, Z => n6891);
   U4565 : NAND2_X1 port map( A1 => n6892, A2 => n6891, ZN => n7007);
   U4566 : XNOR2_X1 port map( A => n7007, B => n6893, ZN => n6900);
   U4567 : NAND2_X1 port map( A1 => n6894, A2 => n6900, ZN => n7066);
   U4568 : INV_X1 port map( A => n6896, ZN => n6897);
   U4569 : XNOR2_X1 port map( A => n4408, B => n6897, ZN => n6899);
   U4570 : XNOR2_X1 port map( A => n6899, B => n7062, ZN => n6902);
   U4571 : INV_X1 port map( A => n6900, ZN => n6901);
   U4572 : NAND2_X1 port map( A1 => n6902, A2 => n6901, ZN => n7067);
   U4573 : NAND2_X1 port map( A1 => n7066, A2 => n7067, ZN => n6907);
   U4574 : INV_X1 port map( A => n6903, ZN => n6904);
   U4575 : XNOR2_X1 port map( A => n6907, B => n8452, ZN => n6908);
   U4576 : NAND2_X1 port map( A1 => n6909, A2 => n6908, ZN => n6987);
   U4577 : NAND2_X1 port map( A1 => n6987, A2 => n6988, ZN => n6928);
   U4578 : NAND2_X1 port map( A1 => n6915, A2 => n8576, ZN => n6912);
   U4579 : NAND2_X1 port map( A1 => n6912, A2 => n6910, ZN => n6914);
   U4580 : NAND2_X1 port map( A1 => n6912, A2 => n8579, ZN => n6913);
   U4581 : OAI211_X1 port map( C1 => n6915, C2 => n8576, A => n6914, B => n6913
                           , ZN => n6924);
   U4582 : XNOR2_X1 port map( A => n8554, B => n6917, ZN => n6938);
   U4583 : INV_X1 port map( A => n6918, ZN => n6937);
   U4584 : XNOR2_X1 port map( A => n6938, B => n6937, ZN => n6975);
   U4585 : NAND2_X1 port map( A1 => n6920, A2 => n6919, ZN => n6922);
   U4587 : NAND2_X1 port map( A1 => n6975, A2 => n6970, ZN => n6923);
   U4588 : NAND2_X1 port map( A1 => n6924, A2 => n6923, ZN => n6985);
   U4589 : INV_X1 port map( A => n6975, ZN => n6926);
   U4590 : NAND2_X1 port map( A1 => n6926, A2 => n6925, ZN => n6990);
   U4591 : NAND2_X1 port map( A1 => n6985, A2 => n6990, ZN => n6927);
   U4592 : XNOR2_X1 port map( A => n6928, B => n6927, ZN => n7364);
   U4593 : NAND2_X1 port map( A1 => n8587, A2 => n8599, ZN => n6930);
   U4594 : OAI211_X1 port map( C1 => n6932, C2 => n6931, A => n6930, B => n6933
                           , ZN => n6936);
   U4595 : INV_X1 port map( A => n8576, ZN => n6934);
   U4596 : XNOR2_X1 port map( A => n6918, B => n6970, ZN => n6939);
   U4598 : XNOR2_X1 port map( A => n6944, B => n6943, ZN => n6974);
   U4599 : NAND2_X1 port map( A1 => n6947, A2 => n8513, ZN => n6966);
   U4600 : INV_X1 port map( A => n6958, ZN => n6955);
   U4601 : OR2_X1 port map( A1 => n6949, A2 => n6948, ZN => n6954);
   U4603 : OAI21_X1 port map( B1 => n8502, B2 => n6951, A => n6950, ZN => n6953
                           );
   U4604 : NAND3_X1 port map( A1 => n6955, A2 => n6954, A3 => n6953, ZN => 
                           n6956);
   U4605 : NAND2_X1 port map( A1 => n6956, A2 => n4421, ZN => n6961);
   U4606 : NAND2_X1 port map( A1 => n6959, A2 => n6958, ZN => n6960);
   U4607 : NAND3_X1 port map( A1 => n6961, A2 => n6957, A3 => n6960, ZN => 
                           n6964);
   U4608 : NAND2_X1 port map( A1 => n6964, A2 => n6963, ZN => n6965);
   U4609 : NAND2_X1 port map( A1 => n6966, A2 => n6965, ZN => n6973);
   U4610 : OAI21_X1 port map( B1 => n6967, B2 => n6945, A => n6973, ZN => n6969
                           );
   U4611 : NAND2_X1 port map( A1 => n6967, A2 => n6945, ZN => n6968);
   U4612 : NAND2_X1 port map( A1 => n6969, A2 => n6968, ZN => n7365);
   U4613 : NAND2_X1 port map( A1 => n7364, A2 => n7365, ZN => n8126);
   U4614 : XNOR2_X1 port map( A => n8598, B => n6970, ZN => n6972);
   U4615 : XNOR2_X1 port map( A => n6973, B => n6972, ZN => n6978);
   U4616 : INV_X1 port map( A => n6974, ZN => n6976);
   U4617 : XNOR2_X1 port map( A => n6976, B => n6975, ZN => n6977);
   U4618 : XNOR2_X1 port map( A => n6978, B => n6977, ZN => n8115);
   U4619 : NAND2_X1 port map( A1 => n6981, A2 => n6979, ZN => n6984);
   U4620 : NAND2_X1 port map( A1 => n6981, A2 => n6980, ZN => n6983);
   U4622 : NAND2_X1 port map( A1 => n8116, A2 => n8115, ZN => n8129);
   U4624 : INV_X1 port map( A => n6987, ZN => n6991);
   U4625 : INV_X1 port map( A => n6985, ZN => n6986);
   U4626 : NAND2_X1 port map( A1 => n6987, A2 => n6986, ZN => n6989);
   U4627 : OAI211_X1 port map( C1 => n6991, C2 => n6990, A => n6989, B => n8464
                           , ZN => n7478);
   U4629 : AOI21_X1 port map( B1 => n6995, B2 => n6994, A => n8473, ZN => n7164
                           );
   U4630 : NAND2_X1 port map( A1 => n6997, A2 => n6996, ZN => n7000);
   U4631 : INV_X1 port map( A => n6998, ZN => n6999);
   U4632 : NAND2_X1 port map( A1 => n7000, A2 => n6999, ZN => n7003);
   U4633 : NAND2_X1 port map( A1 => n7001, A2 => n4435, ZN => n7002);
   U4634 : NAND2_X1 port map( A1 => n7003, A2 => n7002, ZN => n7114);
   U4635 : NAND2_X1 port map( A1 => n7005, A2 => n7004, ZN => n7009);
   U4636 : NAND2_X1 port map( A1 => n7007, A2 => n7006, ZN => n7008);
   U4638 : XNOR2_X1 port map( A => n7114, B => n4465, ZN => n7019);
   U4639 : MUX2_X1 port map( A => n7231, B => n7010, S => n205, Z => n7011);
   U4640 : NAND2_X1 port map( A1 => n7232, A2 => n357, ZN => n7013);
   U4641 : AND2_X1 port map( A1 => n8504, A2 => n8351, ZN => n7128);
   U4642 : NAND2_X1 port map( A1 => n7015, A2 => n7128, ZN => n7147);
   U4643 : NAND2_X1 port map( A1 => n7147, A2 => n7146, ZN => n7018);
   U4644 : MUX2_X1 port map( A => n8476, B => n7559, S => n360, Z => n7017);
   U4645 : MUX2_X1 port map( A => n7227, B => n7439, S => n377, Z => n7016);
   U4646 : NAND2_X1 port map( A1 => n7017, A2 => n7016, ZN => n7144);
   U4647 : XNOR2_X1 port map( A => n7018, B => n7144, ZN => n7115);
   U4648 : XNOR2_X1 port map( A => n7019, B => n8603, ZN => n7074);
   U4649 : INV_X1 port map( A => n7020, ZN => n7028);
   U4650 : INV_X1 port map( A => n7022, ZN => n7024);
   U4651 : AOI21_X1 port map( B1 => n7021, B2 => n7024, A => n4486, ZN => n7026
                           );
   U4652 : NOR2_X1 port map( A1 => n7021, A2 => n7024, ZN => n7025);
   U4653 : OAI22_X1 port map( A1 => n7028, A2 => n7027, B1 => n7026, B2 => 
                           n7025, ZN => n7031);
   U4655 : NAND2_X1 port map( A1 => n7027, A2 => n7028, ZN => n7030);
   U4656 : NAND2_X1 port map( A1 => n7031, A2 => n7030, ZN => n7075);
   U4657 : XNOR2_X1 port map( A => n7074, B => n7075, ZN => n7160);
   U4658 : XNOR2_X1 port map( A => n7164, B => n7160, ZN => n7070);
   U4659 : MUX2_X1 port map( A => n7692, B => n7254, S => n8392, Z => n7032);
   U4660 : NAND2_X1 port map( A1 => n7499, A2 => n4381, ZN => n7033);
   U4662 : MUX2_X1 port map( A => n6460, B => n5226, S => n371, Z => n7036);
   U4663 : NAND2_X1 port map( A1 => n7038, A2 => n7039, ZN => n7108);
   U4664 : INV_X1 port map( A => n7038, ZN => n7041);
   U4665 : INV_X1 port map( A => n7039, ZN => n7040);
   U4666 : NAND2_X1 port map( A1 => n7041, A2 => n7040, ZN => n7110);
   U4667 : NAND2_X1 port map( A1 => n7108, A2 => n7110, ZN => n7046);
   U4668 : NAND2_X1 port map( A1 => n7043, A2 => n7042, ZN => n7045);
   U4669 : NAND2_X1 port map( A1 => n7045, A2 => n7044, ZN => n7109);
   U4670 : XNOR2_X1 port map( A => n7046, B => n7109, ZN => n7059);
   U4671 : MUX2_X1 port map( A => n7086, B => n7047, S => n359, Z => n7049);
   U4672 : MUX2_X1 port map( A => n8559, B => n8582, S => n356, Z => n7048);
   U4673 : NAND2_X1 port map( A1 => n7049, A2 => n7048, ZN => n7134);
   U4674 : INV_X1 port map( A => n7134, ZN => n7137);
   U4675 : MUX2_X1 port map( A => n8469, B => n8596, S => n7506, Z => n7052);
   U4676 : NAND2_X1 port map( A1 => n7052, A2 => n7051, ZN => n7135);
   U4677 : XNOR2_X1 port map( A => n7134, B => n7135, ZN => n7057);
   U4678 : MUX2_X1 port map( A => n8501, B => n7053, S => n363, Z => n7056);
   U4679 : MUX2_X1 port map( A => n4462, B => n7054, S => n8330, Z => n7055);
   U4680 : NAND2_X1 port map( A1 => n7056, A2 => n7055, ZN => n7133);
   U4681 : XNOR2_X1 port map( A => n7133, B => n7057, ZN => n7058);
   U4682 : NAND2_X1 port map( A1 => n7059, A2 => n7058, ZN => n7155);
   U4683 : NAND2_X1 port map( A1 => n7155, A2 => n7156, ZN => n7063);
   U4684 : XNOR2_X1 port map( A => n7063, B => n7153, ZN => n7165);
   U4685 : INV_X1 port map( A => n7064, ZN => n7065);
   U4686 : NAND2_X1 port map( A1 => n7066, A2 => n7065, ZN => n7068);
   U4687 : NAND2_X1 port map( A1 => n7068, A2 => n7067, ZN => n7161);
   U4688 : XNOR2_X1 port map( A => n7167, B => n8602, ZN => n7069);
   U4689 : XNOR2_X1 port map( A => n7070, B => n7069, ZN => n7477);
   U4692 : NAND2_X1 port map( A1 => n8485, A2 => n8456, ZN => n7073);
   U4693 : NAND2_X1 port map( A1 => n7161, A2 => n7073, ZN => n7077);
   U4694 : NAND2_X1 port map( A1 => n8550, A2 => n7075, ZN => n7076);
   U4695 : NAND2_X1 port map( A1 => n7077, A2 => n7076, ZN => n7284);
   U4696 : MUX2_X1 port map( A => n7253, B => n7771, S => n356, Z => n7079);
   U4697 : MUX2_X1 port map( A => n7692, B => n7773, S => n4381, Z => n7078);
   U4698 : NAND2_X1 port map( A1 => n7079, A2 => n7078, ZN => n7237);
   U4699 : MUX2_X1 port map( A => n7195, B => n7080, S => n205, Z => n7082);
   U4700 : MUX2_X1 port map( A => n7324, B => n8465, S => n8349, Z => n7081);
   U4701 : NAND2_X1 port map( A1 => n7082, A2 => n7081, ZN => n7239);
   U4702 : NAND2_X1 port map( A1 => n7051, A2 => n8596, ZN => n7235);
   U4703 : INV_X1 port map( A => n7086, ZN => n7211);
   U4704 : NAND2_X1 port map( A1 => n7211, A2 => n8332, ZN => n7089);
   U4705 : NAND2_X1 port map( A1 => n7089, A2 => n7088, ZN => n7092);
   U4706 : INV_X1 port map( A => n8559, ZN => n7212);
   U4707 : MUX2_X1 port map( A => n7212, B => n7751, S => n359, Z => n7091);
   U4708 : NOR2_X1 port map( A1 => n7092, A2 => n7091, ZN => n7100);
   U4709 : MUX2_X1 port map( A => n7094, B => n7093, S => n372, Z => n7098);
   U4710 : MUX2_X1 port map( A => n7096, B => n7095, S => n360, Z => n7097);
   U4711 : NOR2_X1 port map( A1 => n7098, A2 => n7097, ZN => n7099);
   U4712 : NAND2_X1 port map( A1 => n7100, A2 => n7099, ZN => n7182);
   U4713 : NAND2_X1 port map( A1 => n7182, A2 => n7180, ZN => n7103);
   U4714 : MUX2_X1 port map( A => n8500, B => n7053, S => n371, Z => n7102);
   U4715 : MUX2_X1 port map( A => n4462, B => n7198, S => n8329, Z => n7101);
   U4716 : AND2_X1 port map( A1 => n7102, A2 => n7101, ZN => n7181);
   U4717 : XNOR2_X1 port map( A => n7103, B => n7181, ZN => n7105);
   U4718 : INV_X1 port map( A => n7104, ZN => n7107);
   U4719 : INV_X1 port map( A => n7105, ZN => n7106);
   U4720 : NAND2_X1 port map( A1 => n7107, A2 => n7106, ZN => n7192);
   U4721 : NAND2_X1 port map( A1 => n7191, A2 => n7192, ZN => n7113);
   U4722 : INV_X1 port map( A => n7108, ZN => n7112);
   U4723 : INV_X1 port map( A => n7109, ZN => n7111);
   U4724 : OAI21_X1 port map( B1 => n7112, B2 => n7111, A => n7110, ZN => n7190
                           );
   U4725 : XNOR2_X1 port map( A => n7113, B => n7190, ZN => n7283);
   U4726 : XNOR2_X1 port map( A => n7284, B => n7283, ZN => n7159);
   U4727 : INV_X1 port map( A => n7114, ZN => n7117);
   U4728 : OAI21_X1 port map( B1 => n7117, B2 => n4465, A => n7115, ZN => n7119
                           );
   U4729 : NAND2_X1 port map( A1 => n7117, A2 => n4465, ZN => n7118);
   U4730 : MUX2_X1 port map( A => n7121, B => n4360, S => n7506, Z => n7125);
   U4731 : MUX2_X1 port map( A => n7123, B => n7122, S => n357, Z => n7124);
   U4732 : NAND2_X1 port map( A1 => n7125, A2 => n7124, ZN => n7129);
   U4733 : INV_X1 port map( A => n7128, ZN => n7127);
   U4734 : NAND2_X1 port map( A1 => n4514, A2 => n8392, ZN => n7126);
   U4735 : NAND2_X1 port map( A1 => n7127, A2 => n7126, ZN => n7130);
   U4736 : NAND2_X1 port map( A1 => n7128, A2 => n8392, ZN => n7172);
   U4737 : INV_X1 port map( A => n7129, ZN => n7132);
   U4738 : NAND2_X1 port map( A1 => n7172, A2 => n7130, ZN => n7131);
   U4739 : AOI22_X1 port map( A1 => n7174, A2 => n7172, B1 => n7132, B2 => 
                           n7131, ZN => n7140);
   U4740 : INV_X1 port map( A => n7133, ZN => n7139);
   U4741 : NAND2_X1 port map( A1 => n7134, A2 => n7135, ZN => n7138);
   U4742 : INV_X1 port map( A => n7135, ZN => n7136);
   U4743 : AOI22_X1 port map( A1 => n7139, A2 => n7138, B1 => n7137, B2 => 
                           n7136, ZN => n7141);
   U4744 : NAND2_X1 port map( A1 => n7140, A2 => n7141, ZN => n7186);
   U4748 : NAND2_X1 port map( A1 => n7186, A2 => n7188, ZN => n7150);
   U4749 : INV_X1 port map( A => n7144, ZN => n7145);
   U4750 : NAND2_X1 port map( A1 => n7146, A2 => n7145, ZN => n7148);
   U4751 : XNOR2_X1 port map( A => n7150, B => n7149, ZN => n7151);
   U4752 : NAND2_X1 port map( A1 => n7152, A2 => n7151, ZN => n7276);
   U4753 : NAND2_X1 port map( A1 => n7276, A2 => n7278, ZN => n7158);
   U4754 : NAND2_X1 port map( A1 => n7155, A2 => n7154, ZN => n7157);
   U4755 : NAND2_X1 port map( A1 => n7157, A2 => n7156, ZN => n7277);
   U4756 : XNOR2_X1 port map( A => n7158, B => n7277, ZN => n7286);
   U4757 : XNOR2_X1 port map( A => n7286, B => n7159, ZN => n7371);
   U4759 : AND2_X1 port map( A1 => n8604, A2 => n7165, ZN => n7163);
   U4760 : XNOR2_X1 port map( A => n7163, B => n7162, ZN => n7171);
   U4761 : INV_X1 port map( A => n7164, ZN => n7170);
   U4762 : INV_X1 port map( A => n8602, ZN => n7169);
   U4763 : XNOR2_X1 port map( A => n7167, B => n7160, ZN => n7168);
   U4764 : AOI22_X1 port map( A1 => n7171, A2 => n7170, B1 => n7169, B2 => 
                           n7168, ZN => n7370);
   U4765 : NAND2_X1 port map( A1 => n7370, A2 => n7371, ZN => n8157);
   U4766 : AND2_X1 port map( A1 => n8149, A2 => n8157, ZN => n7480);
   U4767 : INV_X1 port map( A => n7172, ZN => n7173);
   U4768 : MUX2_X1 port map( A => n7253, B => n7771, S => n359, Z => n7176);
   U4769 : MUX2_X1 port map( A => n7692, B => n7773, S => n8326, Z => n7175);
   U4770 : AND2_X1 port map( A1 => n7176, A2 => n7175, ZN => n7178);
   U4771 : NAND2_X1 port map( A1 => n7177, A2 => n7178, ZN => n7264);
   U4772 : INV_X1 port map( A => n7178, ZN => n7179);
   U4773 : NAND2_X1 port map( A1 => n4442, A2 => n7179, ZN => n7263);
   U4774 : NAND2_X1 port map( A1 => n7264, A2 => n7263, ZN => n7184);
   U4775 : NAND2_X1 port map( A1 => n7181, A2 => n7180, ZN => n7183);
   U4776 : AND2_X1 port map( A1 => n7183, A2 => n7182, ZN => n7265);
   U4777 : NAND2_X1 port map( A1 => n7186, A2 => n7185, ZN => n7187);
   U4778 : INV_X1 port map( A => n7355, ZN => n7189);
   U4779 : NAND2_X1 port map( A1 => n7191, A2 => n7190, ZN => n7193);
   U4780 : NAND2_X1 port map( A1 => n7193, A2 => n7192, ZN => n7271);
   U4781 : OAI22_X1 port map( A1 => n7194, A2 => n7271, B1 => n7189, B2 => 
                           n4443, ZN => n7226);
   U4782 : MUX2_X1 port map( A => n7195, B => n4437, S => n7769, Z => n7197);
   U4783 : MUX2_X1 port map( A => n7324, B => n8465, S => n8331, Z => n7196);
   U4784 : NAND2_X1 port map( A1 => n7197, A2 => n7196, ZN => n7341);
   U4785 : XNOR2_X1 port map( A => n7341, B => n7230, ZN => n7201);
   U4786 : MUX2_X1 port map( A => n8500, B => n7053, S => n205, Z => n7200);
   U4787 : MUX2_X1 port map( A => n4462, B => n7198, S => n8349, Z => n7199);
   U4788 : NAND2_X1 port map( A1 => n7200, A2 => n7199, ZN => n7339);
   U4789 : XNOR2_X1 port map( A => n7201, B => n7339, ZN => n7205);
   U4790 : MUX2_X1 port map( A => n8476, B => n7559, S => n371, Z => n7203);
   U4791 : MUX2_X1 port map( A => n7227, B => n7439, S => n363, Z => n7202);
   U4792 : NAND2_X1 port map( A1 => n7203, A2 => n7202, ZN => n7333);
   U4793 : AND2_X1 port map( A1 => n4514, A2 => n8326, ZN => n7334);
   U4794 : NAND2_X1 port map( A1 => n8504, A2 => n4381, ZN => n7330);
   U4795 : XNOR2_X1 port map( A => n7334, B => n7330, ZN => n7204);
   U4796 : XNOR2_X1 port map( A => n7333, B => n7204, ZN => n7206);
   U4797 : NAND2_X1 port map( A1 => n7205, A2 => n7206, ZN => n7320);
   U4798 : NAND2_X1 port map( A1 => n7320, A2 => n7319, ZN => n7225);
   U4799 : MUX2_X1 port map( A => n8500, B => n7053, S => n8423, Z => n7210);
   U4800 : MUX2_X1 port map( A => n4462, B => n7198, S => n8325, Z => n7209);
   U4801 : NAND2_X1 port map( A1 => n7210, A2 => n7209, ZN => n7245);
   U4802 : INV_X1 port map( A => n7245, ZN => n7221);
   U4803 : MUX2_X1 port map( A => n7211, B => n7087, S => n360, Z => n7214);
   U4804 : MUX2_X1 port map( A => n7212, B => n7751, S => n377, Z => n7213);
   U4805 : NOR2_X1 port map( A1 => n7214, A2 => n7213, ZN => n7223);
   U4806 : INV_X1 port map( A => n7223, ZN => n7220);
   U4807 : MUX2_X1 port map( A => n7216, B => n7215, S => n357, Z => n7218);
   U4808 : MUX2_X1 port map( A => n6460, B => n5226, S => n205, Z => n7217);
   U4809 : NOR2_X1 port map( A1 => n7218, A2 => n7217, ZN => n7222);
   U4810 : INV_X1 port map( A => n7222, ZN => n7219);
   U4811 : NAND2_X1 port map( A1 => n7220, A2 => n7219, ZN => n7243);
   U4812 : NAND2_X1 port map( A1 => n7221, A2 => n7243, ZN => n7224);
   U4813 : NAND2_X1 port map( A1 => n7223, A2 => n7222, ZN => n7244);
   U4814 : AND2_X1 port map( A1 => n7224, A2 => n7244, ZN => n7317);
   U4815 : XNOR2_X1 port map( A => n7225, B => n7317, ZN => n7354);
   U4816 : XNOR2_X1 port map( A => n7226, B => n7354, ZN => n7268);
   U4817 : MUX2_X1 port map( A => n8476, B => n7559, S => n363, Z => n7229);
   U4818 : MUX2_X1 port map( A => n7227, B => n7439, S => n372, Z => n7228);
   U4819 : NAND2_X1 port map( A1 => n7229, A2 => n7228, ZN => n7251);
   U4820 : XNOR2_X1 port map( A => n7251, B => n7330, ZN => n7234);
   U4821 : INV_X1 port map( A => n7230, ZN => n7340);
   U4822 : NOR2_X1 port map( A1 => n7232, A2 => n7231, ZN => n7233);
   U4823 : MUX2_X1 port map( A => n7340, B => n7233, S => n8336, Z => n7250);
   U4824 : XNOR2_X1 port map( A => n7234, B => n7250, ZN => n7269);
   U4825 : INV_X1 port map( A => n7235, ZN => n7238);
   U4826 : NAND2_X1 port map( A1 => n7237, A2 => n7236, ZN => n7241);
   U4827 : NAND2_X1 port map( A1 => n7239, A2 => n7238, ZN => n7240);
   U4828 : NAND2_X1 port map( A1 => n7241, A2 => n7240, ZN => n7291);
   U4829 : INV_X1 port map( A => n7291, ZN => n7242);
   U4830 : NAND2_X1 port map( A1 => n7244, A2 => n7243, ZN => n7246);
   U4831 : XNOR2_X1 port map( A => n7246, B => n7245, ZN => n7270);
   U4832 : NAND2_X1 port map( A1 => n7269, A2 => n7242, ZN => n7247);
   U4833 : OAI21_X1 port map( B1 => n7248, B2 => n7270, A => n7247, ZN => n7262
                           );
   U4834 : INV_X1 port map( A => n7250, ZN => n7249);
   U4835 : NAND2_X1 port map( A1 => n7249, A2 => n7330, ZN => n7307);
   U4836 : INV_X1 port map( A => n7330, ZN => n7332);
   U4837 : NAND2_X1 port map( A1 => n7250, A2 => n7332, ZN => n7252);
   U4838 : NAND2_X1 port map( A1 => n7252, A2 => n7251, ZN => n7308);
   U4839 : NAND2_X1 port map( A1 => n7307, A2 => n7308, ZN => n7260);
   U4841 : MUX2_X1 port map( A => n7499, B => n7690, S => n377, Z => n7256);
   U4842 : INV_X1 port map( A => n7254, ZN => n7748);
   U4843 : MUX2_X1 port map( A => n5746, B => n7748, S => n8394, Z => n7255);
   U4844 : NOR2_X1 port map( A1 => n7256, A2 => n7255, ZN => n7309);
   U4845 : MUX2_X1 port map( A => n7665, B => n7556, S => n372, Z => n7258);
   U4846 : MUX2_X1 port map( A => n7696, B => n7695, S => n360, Z => n7257);
   U4847 : NAND2_X1 port map( A1 => n7258, A2 => n7257, ZN => n7306);
   U4848 : XNOR2_X1 port map( A => n7309, B => n7306, ZN => n7259);
   U4849 : XNOR2_X1 port map( A => n7260, B => n7259, ZN => n7261);
   U4850 : NAND2_X1 port map( A1 => n7262, A2 => n7261, ZN => n7351);
   U4851 : NAND2_X1 port map( A1 => n7350, A2 => n7351, ZN => n7267);
   U4852 : INV_X1 port map( A => n7263, ZN => n7266);
   U4853 : OAI21_X1 port map( B1 => n7266, B2 => n7265, A => n7264, ZN => n7349
                           );
   U4855 : XNOR2_X1 port map( A => n7268, B => n4467, ZN => n7378);
   U4856 : OR2_X1 port map( A1 => n7271, A2 => n4443, ZN => n7357);
   U4857 : NAND2_X1 port map( A1 => n7271, A2 => n4443, ZN => n7356);
   U4858 : NAND2_X1 port map( A1 => n7357, A2 => n7356, ZN => n7290);
   U4859 : XNOR2_X1 port map( A => n7290, B => n7355, ZN => n7282);
   U4860 : XNOR2_X1 port map( A => n7270, B => n7269, ZN => n7292);
   U4861 : XNOR2_X1 port map( A => n7292, B => n7242, ZN => n7274);
   U4862 : INV_X1 port map( A => n7274, ZN => n7281);
   U4863 : XNOR2_X1 port map( A => n4443, B => n7355, ZN => n7273);
   U4864 : INV_X1 port map( A => n7271, ZN => n7272);
   U4865 : XNOR2_X1 port map( A => n7273, B => n7272, ZN => n7275);
   U4866 : NAND2_X1 port map( A1 => n7275, A2 => n7274, ZN => n7280);
   U4867 : NAND2_X1 port map( A1 => n7277, A2 => n7276, ZN => n7279);
   U4868 : NAND2_X1 port map( A1 => n7279, A2 => n7278, ZN => n7289);
   U4869 : NAND2_X1 port map( A1 => n7607, A2 => n7378, ZN => n7377);
   U4870 : INV_X1 port map( A => n7283, ZN => n7285);
   U4871 : OAI21_X1 port map( B1 => n7286, B2 => n7285, A => n7284, ZN => n7288
                           );
   U4872 : XNOR2_X1 port map( A => n7290, B => n7289, ZN => n7295);
   U4873 : XNOR2_X1 port map( A => n7355, B => n7291, ZN => n7293);
   U4874 : XNOR2_X1 port map( A => n7293, B => n7292, ZN => n7294);
   U4875 : XNOR2_X1 port map( A => n7295, B => n7294, ZN => n7374);
   U4876 : NOR2_X1 port map( A1 => n7374, A2 => n7373, ZN => n7605);
   U4878 : MUX2_X1 port map( A => n7499, B => n7690, S => n360, Z => n7298);
   U4879 : MUX2_X1 port map( A => n5746, B => n7748, S => n8332, Z => n7297);
   U4880 : MUX2_X1 port map( A => n7665, B => n7556, S => n363, Z => n7300);
   U4881 : MUX2_X1 port map( A => n7696, B => n7695, S => n372, Z => n7299);
   U4882 : AND2_X1 port map( A1 => n7300, A2 => n7299, ZN => n7301);
   U4883 : NAND2_X1 port map( A1 => n7302, A2 => n7301, ZN => n7398);
   U4884 : NAND2_X1 port map( A1 => n7401, A2 => n7398, ZN => n7305);
   U4885 : MUX2_X1 port map( A => n8501, B => n7053, S => n357, Z => n7304);
   U4886 : MUX2_X1 port map( A => n4462, B => n7198, S => n8334, Z => n7303);
   U4887 : AND2_X1 port map( A1 => n7304, A2 => n7303, ZN => n7400);
   U4888 : XNOR2_X1 port map( A => n7305, B => n7400, ZN => n7316);
   U4889 : INV_X1 port map( A => n7316, ZN => n7314);
   U4890 : INV_X1 port map( A => n7306, ZN => n7310);
   U4891 : OAI211_X1 port map( C1 => n7310, C2 => n7309, A => n7308, B => n7307
                           , ZN => n7312);
   U4892 : NAND2_X1 port map( A1 => n7310, A2 => n7309, ZN => n7311);
   U4893 : NAND2_X1 port map( A1 => n7312, A2 => n7311, ZN => n7315);
   U4894 : INV_X1 port map( A => n7315, ZN => n7313);
   U4895 : NAND2_X1 port map( A1 => n7314, A2 => n7313, ZN => n7424);
   U4896 : NAND2_X1 port map( A1 => n7316, A2 => n7315, ZN => n7426);
   U4897 : NAND2_X1 port map( A1 => n7424, A2 => n7426, ZN => n7322);
   U4898 : INV_X1 port map( A => n7317, ZN => n7318);
   U4899 : NAND2_X1 port map( A1 => n7319, A2 => n7318, ZN => n7321);
   U4900 : NAND2_X1 port map( A1 => n7321, A2 => n7320, ZN => n7425);
   U4901 : XNOR2_X1 port map( A => n7322, B => n7425, ZN => n7345);
   U4902 : MUX2_X1 port map( A => n7324, B => n8465, S => n8336, Z => n7326);
   U4903 : NAND2_X1 port map( A1 => n7326, A2 => n7325, ZN => n7389);
   U4904 : NAND2_X1 port map( A1 => n4514, A2 => n8394, ZN => n7466);
   U4905 : XNOR2_X1 port map( A => n7389, B => n7466, ZN => n7329);
   U4906 : MUX2_X1 port map( A => n8476, B => n7559, S => n8423, Z => n7328);
   U4907 : MUX2_X1 port map( A => n7227, B => n7439, S => n371, Z => n7327);
   U4908 : NAND2_X1 port map( A1 => n7328, A2 => n7327, ZN => n7391);
   U4909 : XNOR2_X1 port map( A => n7329, B => n7391, ZN => n7405);
   U4910 : INV_X1 port map( A => n7333, ZN => n7331);
   U4911 : NAND2_X1 port map( A1 => n7331, A2 => n7330, ZN => n7338);
   U4912 : NAND2_X1 port map( A1 => n7333, A2 => n7332, ZN => n7336);
   U4913 : INV_X1 port map( A => n7334, ZN => n7335);
   U4914 : NAND2_X1 port map( A1 => n7336, A2 => n7335, ZN => n7337);
   U4915 : NAND2_X1 port map( A1 => n7338, A2 => n7337, ZN => n7403);
   U4916 : OAI21_X1 port map( B1 => n7340, B2 => n7341, A => n7339, ZN => n7343
                           );
   U4917 : NAND2_X1 port map( A1 => n7341, A2 => n7340, ZN => n7342);
   U4918 : NAND2_X1 port map( A1 => n7343, A2 => n7342, ZN => n7404);
   U4919 : XNOR2_X1 port map( A => n7403, B => n7404, ZN => n7344);
   U4920 : XNOR2_X1 port map( A => n7405, B => n7344, ZN => n7346);
   U4921 : NAND2_X1 port map( A1 => n7345, A2 => n7346, ZN => n7387);
   U4922 : INV_X1 port map( A => n7345, ZN => n7348);
   U4923 : INV_X1 port map( A => n7346, ZN => n7347);
   U4924 : NAND2_X1 port map( A1 => n7348, A2 => n7347, ZN => n7384);
   U4925 : NAND2_X1 port map( A1 => n7387, A2 => n7384, ZN => n7353);
   U4926 : NAND2_X1 port map( A1 => n7350, A2 => n7349, ZN => n7352);
   U4927 : AND2_X1 port map( A1 => n7352, A2 => n7351, ZN => n7385);
   U4928 : INV_X1 port map( A => n7354, ZN => n7360);
   U4929 : NAND2_X1 port map( A1 => n7356, A2 => n7355, ZN => n7358);
   U4930 : NAND2_X1 port map( A1 => n7358, A2 => n7357, ZN => n7359);
   U4931 : OAI21_X1 port map( B1 => n8592, B2 => n7360, A => n7359, ZN => n7363
                           );
   U4932 : NAND2_X1 port map( A1 => n8592, A2 => n7360, ZN => n7362);
   U4933 : AND2_X1 port map( A1 => n7363, A2 => n7362, ZN => n8180);
   U4934 : NAND2_X1 port map( A1 => n8181, A2 => n8180, ZN => n7636);
   U4935 : INV_X1 port map( A => n8555, ZN => n7367);
   U4936 : INV_X1 port map( A => n7365, ZN => n7366);
   U4937 : NAND4_X1 port map( A1 => n7479, A2 => n7480, A3 => n7636, A4 => 
                           n7601, ZN => n7491);
   U4939 : NAND2_X1 port map( A1 => n8541, A2 => n7602, ZN => n7493);
   U4940 : OAI211_X1 port map( C1 => n8111, C2 => n8526, A => n7493, B => n4417
                           , ZN => n7640);
   U4941 : INV_X1 port map( A => n7597, ZN => n7372);
   U4942 : NAND2_X1 port map( A1 => n8585, A2 => n7372, ZN => n7383);
   U4943 : INV_X1 port map( A => n7373, ZN => n7376);
   U4944 : INV_X1 port map( A => n7374, ZN => n7375);
   U4946 : NAND2_X1 port map( A1 => n8168, A2 => n7377, ZN => n7382);
   U4947 : INV_X1 port map( A => n7378, ZN => n7380);
   U4948 : INV_X1 port map( A => n7607, ZN => n7379);
   U4949 : NAND2_X1 port map( A1 => n7380, A2 => n7379, ZN => n8175);
   U4950 : NAND3_X1 port map( A1 => n7383, A2 => n7382, A3 => n7381, ZN => 
                           n7635);
   U4951 : INV_X1 port map( A => n7385, ZN => n7386);
   U4952 : NAND2_X1 port map( A1 => n7384, A2 => n7386, ZN => n7388);
   U4953 : NAND2_X1 port map( A1 => n7388, A2 => n7387, ZN => n7497);
   U4954 : AND2_X1 port map( A1 => n7389, A2 => n7466, ZN => n7390);
   U4955 : OAI22_X1 port map( A1 => n7391, A2 => n7390, B1 => n7466, B2 => 
                           n7389, ZN => n7396);
   U4956 : INV_X1 port map( A => n7771, ZN => n7747);
   U4957 : MUX2_X1 port map( A => n8528, B => n7747, S => n372, Z => n7394);
   U4958 : MUX2_X1 port map( A => n5746, B => n7748, S => n8337, Z => n7393);
   U4959 : NOR2_X1 port map( A1 => n7394, A2 => n7393, ZN => n7395);
   U4960 : NOR2_X1 port map( A1 => n7396, A2 => n7395, ZN => n7453);
   U4961 : INV_X1 port map( A => n7453, ZN => n7397);
   U4962 : NAND2_X1 port map( A1 => n7396, A2 => n7395, ZN => n7452);
   U4963 : NAND2_X1 port map( A1 => n7397, A2 => n7452, ZN => n7402);
   U4964 : INV_X1 port map( A => n7398, ZN => n7399);
   U4965 : AOI21_X1 port map( B1 => n7401, B2 => n7400, A => n7399, ZN => n7454
                           );
   U4966 : XOR2_X1 port map( A => n7402, B => n7454, Z => n7423);
   U4967 : INV_X1 port map( A => n7423, ZN => n7420);
   U4968 : INV_X1 port map( A => n7403, ZN => n7406);
   U4969 : OAI21_X1 port map( B1 => n7406, B2 => n7405, A => n7404, ZN => n7408
                           );
   U4970 : NAND2_X1 port map( A1 => n7406, A2 => n7405, ZN => n7407);
   U4971 : NAND2_X1 port map( A1 => n7408, A2 => n7407, ZN => n7456);
   U4972 : MUX2_X1 port map( A => n8476, B => n7559, S => n205, Z => n7410);
   U4973 : MUX2_X1 port map( A => n8568, B => n7439, S => n8423, Z => n7409);
   U4974 : NAND2_X1 port map( A1 => n7410, A2 => n7409, ZN => n7469);
   U4975 : INV_X1 port map( A => n7466, ZN => n7411);
   U4976 : NAND2_X1 port map( A1 => n8504, A2 => n8332, ZN => n7465);
   U4977 : XNOR2_X1 port map( A => n7411, B => n7465, ZN => n7412);
   U4978 : XNOR2_X1 port map( A => n7469, B => n7412, ZN => n7458);
   U4979 : XNOR2_X1 port map( A => n7456, B => n7458, ZN => n7419);
   U4980 : MUX2_X1 port map( A => n7665, B => n7556, S => n371, Z => n7414);
   U4981 : MUX2_X1 port map( A => n7696, B => n7695, S => n363, Z => n7413);
   U4982 : NAND2_X1 port map( A1 => n7414, A2 => n7413, ZN => n7447);
   U4983 : XNOR2_X1 port map( A => n7447, B => n7444, ZN => n7418);
   U4984 : MUX2_X1 port map( A => n8500, B => n7053, S => n7506, Z => n7417);
   U4985 : MUX2_X1 port map( A => n4462, B => n7198, S => n8331, Z => n7416);
   U4986 : NAND2_X1 port map( A1 => n7417, A2 => n7416, ZN => n7445);
   U4987 : XNOR2_X1 port map( A => n7418, B => n7445, ZN => n7457);
   U4988 : XNOR2_X1 port map( A => n7419, B => n7457, ZN => n7421);
   U4989 : NAND2_X1 port map( A1 => n7420, A2 => n7421, ZN => n7430);
   U4990 : INV_X1 port map( A => n7421, ZN => n7422);
   U4991 : NAND2_X1 port map( A1 => n7423, A2 => n7422, ZN => n7432);
   U4992 : NAND2_X1 port map( A1 => n7430, A2 => n7432, ZN => n7429);
   U4993 : INV_X1 port map( A => n7424, ZN => n7428);
   U4994 : INV_X1 port map( A => n7425, ZN => n7427);
   U4995 : OAI21_X1 port map( B1 => n7428, B2 => n7427, A => n7426, ZN => n7431
                           );
   U4996 : XNOR2_X1 port map( A => n7429, B => n7431, ZN => n7496);
   U4997 : NAND2_X1 port map( A1 => n7497, A2 => n7496, ZN => n7638);
   U4998 : INV_X1 port map( A => n7430, ZN => n7434);
   U4999 : INV_X1 port map( A => n7431, ZN => n7433);
   U5000 : OAI21_X1 port map( B1 => n7434, B2 => n7433, A => n7432, ZN => n7952
                           );
   U5001 : MUX2_X1 port map( A => n4462, B => n7198, S => n8336, Z => n7435);
   U5002 : AND2_X1 port map( A1 => n7053, A2 => n7435, ZN => n7437);
   U5003 : NAND2_X1 port map( A1 => n4514, A2 => n8337, ZN => n7513);
   U5004 : INV_X1 port map( A => n7513, ZN => n7436);
   U5005 : NAND2_X1 port map( A1 => n7437, A2 => n7436, ZN => n7521);
   U5006 : INV_X1 port map( A => n7437, ZN => n7438);
   U5007 : NAND2_X1 port map( A1 => n7438, A2 => n7513, ZN => n7522);
   U5008 : NAND2_X1 port map( A1 => n7521, A2 => n7522, ZN => n7443);
   U5009 : MUX2_X1 port map( A => n8476, B => n7559, S => n357, Z => n7441);
   U5010 : MUX2_X1 port map( A => n8568, B => n7439, S => n205, Z => n7440);
   U5011 : NAND2_X1 port map( A1 => n7441, A2 => n7440, ZN => n7520);
   U5012 : INV_X1 port map( A => n7520, ZN => n7442);
   U5013 : XNOR2_X1 port map( A => n7443, B => n7442, ZN => n7451);
   U5014 : INV_X1 port map( A => n7444, ZN => n7446);
   U5015 : AOI21_X1 port map( B1 => n7447, B2 => n7446, A => n7445, ZN => n7449
                           );
   U5016 : NOR2_X1 port map( A1 => n7447, A2 => n7446, ZN => n7448);
   U5017 : OR2_X1 port map( A1 => n7449, A2 => n7448, ZN => n7450);
   U5018 : OR2_X1 port map( A1 => n7451, A2 => n7450, ZN => n7534);
   U5019 : NAND2_X1 port map( A1 => n7451, A2 => n7450, ZN => n7532);
   U5020 : NAND2_X1 port map( A1 => n7534, A2 => n7532, ZN => n7455);
   U5021 : OAI21_X1 port map( B1 => n7454, B2 => n7453, A => n7452, ZN => n7535
                           );
   U5022 : XNOR2_X1 port map( A => n7455, B => n7535, ZN => n7579);
   U5023 : INV_X1 port map( A => n7456, ZN => n7459);
   U5024 : AOI22_X1 port map( A1 => n7460, A2 => n7459, B1 => n7458, B2 => 
                           n7457, ZN => n7471);
   U5025 : MUX2_X1 port map( A => n8528, B => n7690, S => n363, Z => n7462);
   U5026 : MUX2_X1 port map( A => n5746, B => n7748, S => n8330, Z => n7461);
   U5027 : NOR2_X1 port map( A1 => n7462, A2 => n7461, ZN => n7526);
   U5028 : MUX2_X1 port map( A => n7665, B => n7556, S => n8423, Z => n7464);
   U5029 : MUX2_X1 port map( A => n7696, B => n7695, S => n371, Z => n7463);
   U5030 : NAND2_X1 port map( A1 => n7464, A2 => n7463, ZN => n7530);
   U5031 : XNOR2_X1 port map( A => n7526, B => n7530, ZN => n7470);
   U5032 : NAND2_X1 port map( A1 => n7466, A2 => n7465, ZN => n7468);
   U5033 : NOR2_X1 port map( A1 => n7466, A2 => n7465, ZN => n7467);
   U5034 : AOI21_X1 port map( B1 => n7469, B2 => n7468, A => n7467, ZN => n7527
                           );
   U5035 : XNOR2_X1 port map( A => n7470, B => n7527, ZN => n7472);
   U5036 : NAND2_X1 port map( A1 => n7471, A2 => n7472, ZN => n7578);
   U5037 : INV_X1 port map( A => n7471, ZN => n7474);
   U5038 : INV_X1 port map( A => n7472, ZN => n7473);
   U5039 : NAND2_X1 port map( A1 => n7474, A2 => n7473, ZN => n7576);
   U5040 : NAND2_X1 port map( A1 => n7578, A2 => n7576, ZN => n7475);
   U5041 : XNOR2_X1 port map( A => n7579, B => n7475, ZN => n7951);
   U5042 : NAND2_X1 port map( A1 => n7952, A2 => n7951, ZN => n7643);
   U5043 : NAND2_X1 port map( A1 => n7638, A2 => n7643, ZN => n7476);
   U5044 : AOI21_X1 port map( B1 => n7635, B2 => n7636, A => n7476, ZN => n7482
                           );
   U5045 : AND2_X1 port map( A1 => n7477, A2 => n4448, ZN => n8162);
   U5046 : AND2_X1 port map( A1 => n7479, A2 => n8162, ZN => n7634);
   U5047 : NAND3_X1 port map( A1 => n7634, A2 => n4500, A3 => n7636, ZN => 
                           n7481);
   U5048 : NAND2_X1 port map( A1 => n7855, A2 => n8484, ZN => n7483);
   U5050 : AND2_X1 port map( A1 => n8098, A2 => n7492, ZN => n7484);
   U5051 : AOI21_X1 port map( B1 => n8074, B2 => n6563, A => n7484, ZN => n7486
                           );
   U5052 : AOI21_X1 port map( B1 => n8484, B2 => n6564, A => n7484, ZN => n7485
                           );
   U5053 : AND2_X1 port map( A1 => n7623, A2 => n7734, ZN => n7489);
   U5054 : INV_X1 port map( A => n8484, ZN => n7488);
   U5056 : NOR2_X1 port map( A1 => n7727, A2 => n7491, ZN => n7494);
   U5057 : NAND2_X1 port map( A1 => n7494, A2 => n8578, ZN => n7721);
   U5058 : INV_X1 port map( A => n7721, ZN => n7495);
   U5060 : AND2_X1 port map( A1 => n8561, A2 => n8229, ZN => n7583);
   U5062 : NOR2_X1 port map( A1 => n7497, A2 => n7496, ZN => n7629);
   U5063 : NOR2_X1 port map( A1 => n7952, A2 => n7951, ZN => n7498);
   U5065 : MUX2_X1 port map( A => n7499, B => n7690, S => n371, Z => n7501);
   U5066 : MUX2_X1 port map( A => n5746, B => n7748, S => n8329, Z => n7500);
   U5067 : NOR2_X1 port map( A1 => n7501, A2 => n7500, ZN => n7538);
   U5068 : INV_X1 port map( A => n7538, ZN => n7543);
   U5069 : NAND2_X1 port map( A1 => n7053, A2 => n4462, ZN => n7541);
   U5070 : XNOR2_X1 port map( A => n7543, B => n7541, ZN => n7505);
   U5071 : MUX2_X1 port map( A => n7665, B => n7556, S => n205, Z => n7504);
   U5072 : MUX2_X1 port map( A => n7696, B => n7695, S => n8423, Z => n7503);
   U5073 : NAND2_X1 port map( A1 => n7504, A2 => n7503, ZN => n7539);
   U5074 : XNOR2_X1 port map( A => n7505, B => n7539, ZN => n7519);
   U5075 : INV_X1 port map( A => n7519, ZN => n7517);
   U5076 : MUX2_X1 port map( A => n8476, B => n7559, S => n7506, Z => n7510);
   U5077 : MUX2_X1 port map( A => n6800, B => n7439, S => n357, Z => n7509);
   U5078 : NAND2_X1 port map( A1 => n7510, A2 => n7509, ZN => n7554);
   U5079 : NAND2_X1 port map( A1 => n4514, A2 => n8330, ZN => n7512);
   U5080 : NOR2_X1 port map( A1 => n7513, A2 => n7512, ZN => n7552);
   U5081 : NAND2_X1 port map( A1 => n7513, A2 => n7512, ZN => n7553);
   U5082 : INV_X1 port map( A => n7553, ZN => n7514);
   U5083 : NOR2_X1 port map( A1 => n7552, A2 => n7514, ZN => n7515);
   U5084 : XNOR2_X1 port map( A => n7554, B => n7515, ZN => n7518);
   U5085 : INV_X1 port map( A => n7518, ZN => n7516);
   U5086 : NAND2_X1 port map( A1 => n7517, A2 => n7516, ZN => n7568);
   U5087 : NAND2_X1 port map( A1 => n7519, A2 => n7518, ZN => n7567);
   U5088 : NAND2_X1 port map( A1 => n7568, A2 => n7567, ZN => n7525);
   U5089 : NAND2_X1 port map( A1 => n7521, A2 => n7520, ZN => n7523);
   U5090 : NAND2_X1 port map( A1 => n7523, A2 => n7522, ZN => n7566);
   U5091 : INV_X1 port map( A => n7566, ZN => n7524);
   U5092 : XNOR2_X1 port map( A => n7525, B => n7524, ZN => n7537);
   U5093 : INV_X1 port map( A => n7527, ZN => n7531);
   U5094 : INV_X1 port map( A => n7530, ZN => n7528);
   U5095 : OAI21_X1 port map( B1 => n7528, B2 => n7527, A => n7526, ZN => n7529
                           );
   U5096 : OAI21_X1 port map( B1 => n7531, B2 => n7530, A => n7529, ZN => n7536
                           );
   U5097 : NOR2_X1 port map( A1 => n7537, A2 => n7536, ZN => n7571);
   U5098 : INV_X1 port map( A => n7532, ZN => n7533);
   U5099 : AOI21_X1 port map( B1 => n7535, B2 => n7534, A => n7533, ZN => n7574
                           );
   U5100 : NAND2_X1 port map( A1 => n7537, A2 => n7536, ZN => n7572);
   U5102 : NAND2_X1 port map( A1 => n7538, A2 => n7541, ZN => n7540);
   U5103 : NAND2_X1 port map( A1 => n7540, A2 => n7539, ZN => n7545);
   U5104 : INV_X1 port map( A => n7541, ZN => n7542);
   U5105 : NAND2_X1 port map( A1 => n7543, A2 => n7542, ZN => n7544);
   U5106 : NAND2_X1 port map( A1 => n7545, A2 => n7544, ZN => n7551);
   U5107 : INV_X1 port map( A => n7551, ZN => n7548);
   U5108 : MUX2_X1 port map( A => n8528, B => n7747, S => n8423, Z => n7547);
   U5109 : MUX2_X1 port map( A => n5746, B => n7748, S => n8325, Z => n7546);
   U5110 : NOR2_X1 port map( A1 => n7547, A2 => n7546, ZN => n7549);
   U5111 : NAND2_X1 port map( A1 => n7548, A2 => n7549, ZN => n7675);
   U5112 : INV_X1 port map( A => n7549, ZN => n7550);
   U5113 : NAND2_X1 port map( A1 => n7551, A2 => n7550, ZN => n7676);
   U5114 : NAND2_X1 port map( A1 => n7675, A2 => n7676, ZN => n7555);
   U5115 : AOI21_X1 port map( B1 => n7554, B2 => n7553, A => n7552, ZN => n7673
                           );
   U5116 : XNOR2_X1 port map( A => n7555, B => n7673, ZN => n7562);
   U5117 : MUX2_X1 port map( A => n7665, B => n7556, S => n357, Z => n7558);
   U5118 : MUX2_X1 port map( A => n7696, B => n7695, S => n205, Z => n7557);
   U5119 : AND2_X1 port map( A1 => n7558, A2 => n7557, ZN => n7663);
   U5120 : AND2_X1 port map( A1 => n4514, A2 => n8329, ZN => n7686);
   U5121 : NAND2_X1 port map( A1 => n7559, A2 => n7227, ZN => n7560);
   U5122 : MUX2_X1 port map( A => n7659, B => n7560, S => n8336, Z => n7561);
   U5123 : INV_X1 port map( A => n7561, ZN => n7662);
   U5124 : NAND2_X1 port map( A1 => n7562, A2 => n7563, ZN => n7653);
   U5125 : INV_X1 port map( A => n7562, ZN => n7565);
   U5126 : INV_X1 port map( A => n7563, ZN => n7564);
   U5127 : NAND2_X1 port map( A1 => n7565, A2 => n7564, ZN => n7654);
   U5128 : NAND2_X1 port map( A1 => n7653, A2 => n7654, ZN => n7570);
   U5129 : NAND2_X1 port map( A1 => n7567, A2 => n7566, ZN => n7569);
   U5130 : NAND2_X1 port map( A1 => n7569, A2 => n7568, ZN => n7652);
   U5131 : XNOR2_X1 port map( A => n7570, B => n7652, ZN => n8205);
   U5132 : XNOR2_X1 port map( A => n7712, B => n8205, ZN => n7587);
   U5133 : INV_X1 port map( A => n7571, ZN => n7573);
   U5134 : NAND2_X1 port map( A1 => n7573, A2 => n7572, ZN => n7575);
   U5135 : XOR2_X1 port map( A => n7575, B => n7574, Z => n7709);
   U5136 : INV_X1 port map( A => n8562, ZN => n7580);
   U5137 : INV_X1 port map( A => n7576, ZN => n7577);
   U5138 : AOI21_X1 port map( B1 => n7579, B2 => n7578, A => n7577, ZN => n7707
                           );
   U5139 : NAND2_X1 port map( A1 => n7580, A2 => n7707, ZN => n8207);
   U5143 : NAND2_X1 port map( A1 => n4414, A2 => n4412, ZN => n7956);
   U5144 : INV_X1 port map( A => n7707, ZN => n7582);
   U5145 : NAND2_X1 port map( A1 => n7709, A2 => n7582, ZN => n8213);
   U5146 : INV_X1 port map( A => n7587, ZN => n7586);
   U5147 : AND2_X1 port map( A1 => n8213, A2 => n7586, ZN => n7589);
   U5148 : NAND3_X1 port map( A1 => n7583, A2 => n7956, A3 => n7589, ZN => 
                           n7592);
   U5150 : NAND3_X1 port map( A1 => n8110, A2 => n8601, A3 => n7585, ZN => 
                           n7591);
   U5151 : INV_X1 port map( A => n8208, ZN => n7633);
   U5152 : OAI22_X1 port map( A1 => n8207, A2 => n7587, B1 => n8213, B2 => 
                           n7586, ZN => n7588);
   U5153 : AOI21_X1 port map( B1 => n7633, B2 => n7589, A => n7588, ZN => n7590
                           );
   U5154 : NAND4_X1 port map( A1 => n8096, A2 => n8146, A3 => n7595, A4 => 
                           n4432, ZN => n8152);
   U5155 : INV_X1 port map( A => n8175, ZN => n7596);
   U5156 : NOR2_X1 port map( A1 => n8168, A2 => n7596, ZN => n7598);
   U5157 : NAND2_X1 port map( A1 => n7598, A2 => n7597, ZN => n7612);
   U5158 : OR2_X1 port map( A1 => n7612, A2 => n8162, ZN => n8186);
   U5159 : INV_X1 port map( A => n7613, ZN => n7600);
   U5161 : INV_X1 port map( A => n7625, ZN => n7617);
   U5162 : INV_X1 port map( A => n4485, ZN => n7604);
   U5163 : INV_X1 port map( A => n7727, ZN => n8099);
   U5165 : INV_X1 port map( A => n8147, ZN => n8127);
   U5166 : NAND3_X1 port map( A1 => n8099, A2 => n8127, A3 => n4485, ZN => 
                           n7603);
   U5167 : OAI211_X1 port map( C1 => n8146, C2 => n7604, A => n7625, B => n7603
                           , ZN => n7616);
   U5168 : OAI21_X1 port map( B1 => n7606, B2 => n7608, A => n7607, ZN => n7610
                           );
   U5169 : NAND2_X1 port map( A1 => n7606, A2 => n7608, ZN => n7609);
   U5170 : AND2_X1 port map( A1 => n7610, A2 => n7609, ZN => n7611);
   U5171 : OAI21_X1 port map( B1 => n7612, B2 => n4500, A => n7611, ZN => n8189
                           );
   U5172 : INV_X1 port map( A => n7636, ZN => n7614);
   U5173 : OAI21_X1 port map( B1 => n8189, B2 => n7614, A => n7613, ZN => n7615
                           );
   U5174 : NOR2_X1 port map( A1 => n7619, A2 => n7618, ZN => n7624);
   U5175 : INV_X1 port map( A => n7620, ZN => n7621);
   U5176 : NAND3_X1 port map( A1 => n8527, A2 => n7624, A3 => n4532, ZN => 
                           n8145);
   U5177 : NAND2_X1 port map( A1 => n4438, A2 => n7625, ZN => n7626);
   U5178 : NAND2_X1 port map( A1 => n4447, A2 => n7737, ZN => n8144);
   U5179 : NAND2_X1 port map( A1 => n7628, A2 => n7627, ZN => n7632);
   U5180 : INV_X1 port map( A => n7638, ZN => n7630);
   U5181 : OR2_X1 port map( A1 => n7630, A2 => n7959, ZN => n7631);
   U5182 : XNOR2_X1 port map( A => n7632, B => n7631, ZN => I2_dtemp_39_port);
   U5183 : AND2_X1 port map( A1 => n8207, A2 => n8213, ZN => n7642);
   U5184 : NAND2_X1 port map( A1 => n4418, A2 => n7956, ZN => n7963);
   U5185 : AND2_X1 port map( A1 => n7634, A2 => n4500, ZN => n7637);
   U5186 : OAI21_X1 port map( B1 => n7637, B2 => n4483, A => n7636, ZN => n7639
                           );
   U5187 : AND3_X1 port map( A1 => n7640, A2 => n7639, A3 => n7638, ZN => n7960
                           );
   U5188 : NAND3_X1 port map( A1 => n7960, A2 => n7642, A3 => n7643, ZN => 
                           n7641);
   U5189 : OR2_X1 port map( A1 => n7963, A2 => n7641, ZN => n7648);
   U5190 : INV_X1 port map( A => n7642, ZN => n7644);
   U5191 : NAND4_X1 port map( A1 => n8605, A2 => n7960, A3 => n7643, A4 => 
                           n7644, ZN => n7646);
   U5192 : XNOR2_X1 port map( A => n8208, B => n7644, ZN => n7645);
   U5193 : NAND2_X1 port map( A1 => n7646, A2 => n7645, ZN => n7647);
   U5194 : AND3_X1 port map( A1 => n7648, A2 => n7649, A3 => n7647, ZN => 
                           I2_dtemp_41_port);
   U5196 : NAND2_X1 port map( A1 => n7653, A2 => n7652, ZN => n7655);
   U5197 : NAND2_X1 port map( A1 => n7655, A2 => n7654, ZN => n7711);
   U5198 : MUX2_X1 port map( A => n7499, B => n7690, S => n205, Z => n7657);
   U5199 : MUX2_X1 port map( A => n5746, B => n7748, S => n8349, Z => n7656);
   U5200 : NOR2_X1 port map( A1 => n7657, A2 => n7656, ZN => n7658);
   U5201 : NAND2_X1 port map( A1 => n7658, A2 => n7659, ZN => n7754);
   U5202 : INV_X1 port map( A => n7658, ZN => n7661);
   U5203 : INV_X1 port map( A => n7659, ZN => n7660);
   U5204 : NAND2_X1 port map( A1 => n7661, A2 => n7660, ZN => n7704);
   U5205 : NAND2_X1 port map( A1 => n7754, A2 => n7704, ZN => n7664);
   U5206 : FA_X1 port map( A => n7663, B => n7686, CI => n7662, CO => n7703, S 
                           => n7563);
   U5207 : XNOR2_X1 port map( A => n7664, B => n7703, ZN => n7669);
   U5208 : MUX2_X1 port map( A => n7665, B => n7556, S => n7769, Z => n7667);
   U5209 : MUX2_X1 port map( A => n7696, B => n7695, S => n357, Z => n7666);
   U5210 : NAND2_X1 port map( A1 => n7667, A2 => n7666, ZN => n7683);
   U5211 : NAND2_X1 port map( A1 => n4514, A2 => n8325, ZN => n7684);
   U5212 : XNOR2_X1 port map( A => n7686, B => n7684, ZN => n7668);
   U5213 : XNOR2_X1 port map( A => n7683, B => n7668, ZN => n7670);
   U5214 : NAND2_X1 port map( A1 => n7669, A2 => n7670, ZN => n7679);
   U5215 : INV_X1 port map( A => n7669, ZN => n7672);
   U5216 : INV_X1 port map( A => n7670, ZN => n7671);
   U5217 : NAND2_X1 port map( A1 => n7672, A2 => n7671, ZN => n7681);
   U5218 : NAND2_X1 port map( A1 => n7679, A2 => n7681, ZN => n7678);
   U5219 : INV_X1 port map( A => n7673, ZN => n7674);
   U5220 : NAND2_X1 port map( A1 => n7675, A2 => n7674, ZN => n7677);
   U5221 : NAND2_X1 port map( A1 => n7677, A2 => n7676, ZN => n7680);
   U5222 : XNOR2_X1 port map( A => n7678, B => n7680, ZN => n8240);
   U5223 : OR2_X1 port map( A1 => n7711, A2 => n8240, ZN => n8232);
   U5224 : NAND2_X1 port map( A1 => n7680, A2 => n7679, ZN => n7682);
   U5225 : NAND2_X1 port map( A1 => n7682, A2 => n7681, ZN => n7714);
   U5226 : INV_X1 port map( A => n7683, ZN => n7689);
   U5227 : INV_X1 port map( A => n7684, ZN => n7685);
   U5228 : NAND2_X1 port map( A1 => n7686, A2 => n7685, ZN => n7688);
   U5229 : NOR2_X1 port map( A1 => n7686, A2 => n7685, ZN => n7687);
   U5230 : AOI21_X1 port map( B1 => n7689, B2 => n7688, A => n7687, ZN => n7700
                           );
   U5231 : MUX2_X1 port map( A => n8528, B => n7690, S => n357, Z => n7691);
   U5232 : INV_X1 port map( A => n7691, ZN => n7694);
   U5233 : MUX2_X1 port map( A => n7692, B => n7773, S => n8334, Z => n7693);
   U5234 : NAND2_X1 port map( A1 => n7694, A2 => n7693, ZN => n7742);
   U5235 : MUX2_X1 port map( A => n7696, B => n7695, S => n7506, Z => n7697);
   U5236 : NAND2_X1 port map( A1 => n7556, A2 => n7697, ZN => n7743);
   U5237 : NAND2_X1 port map( A1 => A_SIG_23_port, A2 => n8349, ZN => n7776);
   U5238 : XNOR2_X1 port map( A => n7743, B => n7776, ZN => n7698);
   U5239 : XNOR2_X1 port map( A => n7742, B => n7698, ZN => n7699);
   U5240 : NAND2_X1 port map( A1 => n7700, A2 => n7699, ZN => n7758);
   U5241 : INV_X1 port map( A => n7699, ZN => n7702);
   U5242 : INV_X1 port map( A => n7700, ZN => n7701);
   U5243 : NAND2_X1 port map( A1 => n7702, A2 => n7701, ZN => n7759);
   U5244 : NAND2_X1 port map( A1 => n7758, A2 => n7759, ZN => n7706);
   U5245 : NAND2_X1 port map( A1 => n7704, A2 => n7703, ZN => n7756);
   U5246 : AND2_X1 port map( A1 => n7756, A2 => n7754, ZN => n7705);
   U5247 : XNOR2_X1 port map( A => n7706, B => n7705, ZN => n7713);
   U5248 : OR2_X1 port map( A1 => n7714, A2 => n7713, ZN => n8231);
   U5249 : AND2_X1 port map( A1 => n8232, A2 => n8231, ZN => n7730);
   U5250 : NAND2_X1 port map( A1 => n7730, A2 => n7707, ZN => n7708);
   U5251 : NOR2_X1 port map( A1 => n8562, A2 => n7708, ZN => n7718);
   U5252 : INV_X1 port map( A => n8205, ZN => n7710);
   U5253 : NAND2_X1 port map( A1 => n7712, A2 => n7710, ZN => n8214);
   U5254 : INV_X1 port map( A => n8231, ZN => n7716);
   U5255 : NAND2_X1 port map( A1 => n7711, A2 => n8240, ZN => n8238);
   U5256 : INV_X1 port map( A => n7712, ZN => n8206);
   U5257 : NAND4_X1 port map( A1 => n8206, A2 => n8205, A3 => n8232, A4 => 
                           n8231, ZN => n7715);
   U5258 : NAND2_X1 port map( A1 => n7714, A2 => n7713, ZN => n8230);
   U5259 : OAI211_X1 port map( C1 => n7716, C2 => n8238, A => n7715, B => n8230
                           , ZN => n7717);
   U5260 : AOI21_X1 port map( B1 => n7718, B2 => n8214, A => n7717, ZN => n7732
                           );
   U5261 : INV_X1 port map( A => n7728, ZN => n7719);
   U5262 : NAND3_X1 port map( A1 => n8590, A2 => n4482, A3 => n7719, ZN => 
                           n7722);
   U5263 : NOR2_X1 port map( A1 => n7722, A2 => n7721, ZN => n7725);
   U5265 : NAND2_X1 port map( A1 => n4417, A2 => n8578, ZN => n8212);
   U5266 : OR2_X1 port map( A1 => n7728, A2 => n7727, ZN => n7729);
   U5268 : NAND3_X1 port map( A1 => n8213, A2 => n7730, A3 => n8214, ZN => 
                           n7731);
   U5269 : NAND2_X1 port map( A1 => n7732, A2 => n7731, ZN => n7988);
   U5271 : INV_X1 port map( A => n8527, ZN => n7740);
   U5272 : AND2_X1 port map( A1 => n7736, A2 => n7735, ZN => n7738);
   U5273 : NAND2_X1 port map( A1 => n7738, A2 => n7737, ZN => n7739);
   U5275 : INV_X1 port map( A => n7742, ZN => n7746);
   U5276 : NOR2_X1 port map( A1 => n7743, A2 => n7776, ZN => n7745);
   U5277 : INV_X1 port map( A => n7743, ZN => n7744);
   U5278 : INV_X1 port map( A => n7776, ZN => n7778);
   U5279 : OAI22_X1 port map( A1 => n7746, A2 => n7745, B1 => n7744, B2 => 
                           n7778, ZN => n7762);
   U5280 : MUX2_X1 port map( A => n8528, B => n7747, S => n7769, Z => n7750);
   U5281 : MUX2_X1 port map( A => n5746, B => n7748, S => n8331, Z => n7749);
   U5282 : NOR2_X1 port map( A1 => n7750, A2 => n7749, ZN => n7763);
   U5283 : XNOR2_X1 port map( A => n7762, B => n7763, ZN => n7753);
   U5284 : OR2_X1 port map( A1 => n7751, A2 => n7087, ZN => n7777);
   U5285 : AND2_X1 port map( A1 => n4514, A2 => n8334, ZN => n7780);
   U5286 : XNOR2_X1 port map( A => n7780, B => n7776, ZN => n7752);
   U5287 : XNOR2_X1 port map( A => n7777, B => n7752, ZN => n7764);
   U5288 : XNOR2_X1 port map( A => n7753, B => n7764, ZN => n7985);
   U5289 : INV_X1 port map( A => n7754, ZN => n7755);
   U5290 : NAND2_X1 port map( A1 => n7758, A2 => n7755, ZN => n7761);
   U5291 : INV_X1 port map( A => n7756, ZN => n7757);
   U5292 : NAND2_X1 port map( A1 => n7758, A2 => n7757, ZN => n7760);
   U5293 : NAND3_X1 port map( A1 => n7761, A2 => n7760, A3 => n7759, ZN => 
                           n7984);
   U5294 : NAND2_X1 port map( A1 => n7985, A2 => n7984, ZN => n7970);
   U5295 : INV_X1 port map( A => n7762, ZN => n7768);
   U5296 : INV_X1 port map( A => n7763, ZN => n7765);
   U5297 : NAND2_X1 port map( A1 => n7765, A2 => n7764, ZN => n7767);
   U5298 : NOR2_X1 port map( A1 => n7765, A2 => n7764, ZN => n7766);
   U5299 : AOI21_X1 port map( B1 => n7768, B2 => n7767, A => n7766, ZN => n7783
                           );
   U5300 : NAND2_X1 port map( A1 => n5746, A2 => n7769, ZN => n7770);
   U5301 : NAND2_X1 port map( A1 => n7771, A2 => n7770, ZN => n7772);
   U5302 : NAND2_X1 port map( A1 => n7772, A2 => n8331, ZN => n7803);
   U5303 : INV_X1 port map( A => n7772, ZN => n7791);
   U5304 : NAND2_X1 port map( A1 => n4514, A2 => n8331, ZN => n7790);
   U5305 : OAI21_X1 port map( B1 => n7773, B2 => n7506, A => n7790, ZN => n7774
                           );
   U5306 : INV_X1 port map( A => n7774, ZN => n7775);
   U5307 : NAND2_X1 port map( A1 => n7791, A2 => n7775, ZN => n7788);
   U5308 : NAND2_X1 port map( A1 => n7803, A2 => n7788, ZN => n7782);
   U5309 : NAND2_X1 port map( A1 => n7777, A2 => n7776, ZN => n7781);
   U5310 : INV_X1 port map( A => n7777, ZN => n7779);
   U5311 : AOI22_X1 port map( A1 => n7781, A2 => n7780, B1 => n7779, B2 => 
                           n7778, ZN => n7797);
   U5312 : XNOR2_X1 port map( A => n7782, B => n7797, ZN => n7784);
   U5313 : AND2_X1 port map( A1 => n7783, A2 => n7784, ZN => n7968);
   U5314 : INV_X1 port map( A => n7783, ZN => n7786);
   U5315 : INV_X1 port map( A => n7784, ZN => n7785);
   U5316 : NAND2_X1 port map( A1 => n7786, A2 => n7785, ZN => n7967);
   U5317 : OAI21_X1 port map( B1 => n7970, B2 => n7968, A => n7967, ZN => n7806
                           );
   U5318 : INV_X1 port map( A => n7806, ZN => n7795);
   U5319 : XNOR2_X1 port map( A => n5748, B => n7769, ZN => n7787);
   U5320 : AND2_X1 port map( A1 => n7787, A2 => n8504, ZN => n7789);
   U5321 : NOR2_X1 port map( A1 => n7788, A2 => n7789, ZN => n7793);
   U5322 : INV_X1 port map( A => n7789, ZN => n7802);
   U5323 : AOI21_X1 port map( B1 => n7791, B2 => n7790, A => n7802, ZN => n7792
                           );
   U5324 : AOI21_X1 port map( B1 => n7793, B2 => n7797, A => n7792, ZN => n7798
                           );
   U5325 : INV_X1 port map( A => n7798, ZN => n7794);
   U5326 : AND2_X1 port map( A1 => n7795, A2 => n7794, ZN => n7796);
   U5327 : AOI21_X1 port map( B1 => n7803, B2 => n7802, A => n7797, ZN => n7799
                           );
   U5328 : NOR2_X1 port map( A1 => n7799, A2 => n7794, ZN => n7805);
   U5329 : INV_X1 port map( A => n7984, ZN => n7973);
   U5330 : INV_X1 port map( A => n7985, ZN => n7976);
   U5331 : NAND2_X1 port map( A1 => n7973, A2 => n7976, ZN => n7971);
   U5332 : INV_X1 port map( A => n7968, ZN => n7800);
   U5333 : NAND3_X1 port map( A1 => n7795, A2 => n7794, A3 => n7801, ZN => 
                           n7808);
   U5334 : NOR2_X1 port map( A1 => n7803, A2 => n7802, ZN => n7804);
   U5335 : AOI21_X1 port map( B1 => n7806, B2 => n7805, A => n7804, ZN => n7807
                           );
   U5336 : NOR2_X1 port map( A1 => FP_B(24), A2 => FP_B(23), ZN => n7812);
   U5337 : NOR2_X1 port map( A1 => FP_B(26), A2 => FP_B(25), ZN => n7811);
   U5338 : NOR2_X1 port map( A1 => FP_B(28), A2 => FP_B(27), ZN => n7810);
   U5339 : NOR2_X1 port map( A1 => FP_B(30), A2 => FP_B(29), ZN => n7809);
   U5340 : NAND4_X1 port map( A1 => n7812, A2 => n7811, A3 => n7810, A4 => 
                           n7809, ZN => I1_I1_N13);
   U5341 : NOR2_X1 port map( A1 => FP_A(24), A2 => FP_A(23), ZN => n7816);
   U5342 : NOR2_X1 port map( A1 => FP_A(26), A2 => FP_A(25), ZN => n7815);
   U5343 : NOR2_X1 port map( A1 => FP_A(28), A2 => FP_A(27), ZN => n7814);
   U5344 : NOR2_X1 port map( A1 => FP_A(30), A2 => FP_A(29), ZN => n7813);
   U5345 : NAND4_X1 port map( A1 => n7816, A2 => n7815, A3 => n7814, A4 => 
                           n7813, ZN => I1_I0_N13);
   U5346 : NOR2_X1 port map( A1 => FP_B(16), A2 => FP_B(15), ZN => n7820);
   U5347 : NOR2_X1 port map( A1 => FP_B(14), A2 => FP_B(13), ZN => n7819);
   U5348 : NOR2_X1 port map( A1 => FP_B(12), A2 => FP_B(11), ZN => n7818);
   U5349 : NOR2_X1 port map( A1 => FP_B(10), A2 => FP_B(9), ZN => n7817);
   U5350 : AND4_X1 port map( A1 => n7820, A2 => n7819, A3 => n7818, A4 => n7817
                           , ZN => n7832);
   U5351 : NOR2_X1 port map( A1 => FP_B(22), A2 => FP_B(21), ZN => n7824);
   U5352 : NOR2_X1 port map( A1 => FP_B(20), A2 => FP_B(19), ZN => n7823);
   U5353 : NOR2_X1 port map( A1 => FP_B(18), A2 => FP_B(17), ZN => n7822);
   U5354 : INV_X1 port map( A => FP_B(0), ZN => n7821);
   U5355 : AND4_X1 port map( A1 => n7824, A2 => n7823, A3 => n7822, A4 => n7821
                           , ZN => n7831);
   U5356 : NOR2_X1 port map( A1 => FP_B(8), A2 => FP_B(7), ZN => n7826);
   U5357 : NOR2_X1 port map( A1 => FP_B(6), A2 => FP_B(5), ZN => n7825);
   U5358 : AND2_X1 port map( A1 => n7826, A2 => n7825, ZN => n7830);
   U5359 : NOR2_X1 port map( A1 => FP_B(4), A2 => FP_B(3), ZN => n7828);
   U5360 : NOR2_X1 port map( A1 => FP_B(2), A2 => FP_B(1), ZN => n7827);
   U5361 : AND2_X1 port map( A1 => n7828, A2 => n7827, ZN => n7829);
   U5362 : NAND4_X1 port map( A1 => n7832, A2 => n7831, A3 => n7830, A4 => 
                           n7829, ZN => n8281);
   U5363 : INV_X1 port map( A => n8281, ZN => n7999);
   U5364 : NAND4_X1 port map( A1 => FP_B(24), A2 => FP_B(23), A3 => FP_B(26), 
                           A4 => FP_B(25), ZN => n7834);
   U5365 : NAND4_X1 port map( A1 => FP_B(28), A2 => FP_B(27), A3 => FP_B(30), 
                           A4 => FP_B(29), ZN => n7833);
   U5366 : NOR2_X1 port map( A1 => n7834, A2 => n7833, ZN => n8280);
   U5367 : NAND2_X1 port map( A1 => n7999, A2 => n8280, ZN => n8283);
   U5368 : INV_X1 port map( A => n8283, ZN => n7852);
   U5369 : NOR2_X1 port map( A1 => FP_A(14), A2 => FP_A(15), ZN => n7838);
   U5370 : NOR2_X1 port map( A1 => FP_A(16), A2 => FP_A(17), ZN => n7837);
   U5371 : NOR2_X1 port map( A1 => FP_A(18), A2 => FP_A(19), ZN => n7836);
   U5372 : NOR2_X1 port map( A1 => FP_A(20), A2 => FP_A(21), ZN => n7835);
   U5373 : AND4_X1 port map( A1 => n7838, A2 => n7837, A3 => n7836, A4 => n7835
                           , ZN => n7848);
   U5374 : NOR2_X1 port map( A1 => FP_A(6), A2 => FP_A(7), ZN => n7842);
   U5375 : NOR2_X1 port map( A1 => FP_A(8), A2 => FP_A(9), ZN => n7841);
   U5376 : NOR2_X1 port map( A1 => FP_A(10), A2 => FP_A(11), ZN => n7840);
   U5377 : NOR2_X1 port map( A1 => FP_A(12), A2 => FP_A(13), ZN => n7839);
   U5378 : AND4_X1 port map( A1 => n7842, A2 => n7841, A3 => n7840, A4 => n7839
                           , ZN => n7847);
   U5379 : NOR3_X1 port map( A1 => FP_A(22), A2 => FP_A(0), A3 => FP_A(1), ZN 
                           => n7846);
   U5380 : NOR2_X1 port map( A1 => FP_A(2), A2 => FP_A(3), ZN => n7844);
   U5381 : NOR2_X1 port map( A1 => FP_A(4), A2 => FP_A(5), ZN => n7843);
   U5382 : AND2_X1 port map( A1 => n7844, A2 => n7843, ZN => n7845);
   U5383 : NAND4_X1 port map( A1 => n7848, A2 => n7847, A3 => n7846, A4 => 
                           n7845, ZN => n8282);
   U5384 : NOR2_X1 port map( A1 => n8282, A2 => I1_I0_N13, ZN => n7997);
   U5385 : NAND4_X1 port map( A1 => FP_A(24), A2 => FP_A(23), A3 => FP_A(26), 
                           A4 => FP_A(25), ZN => n7850);
   U5386 : NAND4_X1 port map( A1 => FP_A(28), A2 => FP_A(27), A3 => FP_A(30), 
                           A4 => FP_A(29), ZN => n7849);
   U5387 : NOR2_X1 port map( A1 => n7850, A2 => n7849, ZN => n8284);
   U5388 : INV_X1 port map( A => n8284, ZN => n7853);
   U5389 : NOR2_X1 port map( A1 => I1_I1_N13, A2 => n7853, ZN => n7851);
   U5390 : AOI22_X1 port map( A1 => n7852, A2 => n7997, B1 => n7999, B2 => 
                           n7851, ZN => n8287);
   U5391 : OAI21_X1 port map( B1 => n8282, B2 => n7853, A => n8283, ZN => n7854
                           );
   U5392 : AND2_X1 port map( A1 => n8287, A2 => n7854, ZN => I1_isINF_int);
   U5393 : INV_X1 port map( A => n8490, ZN => n7856);
   U5394 : NOR2_X1 port map( A1 => n7856, A2 => n8575, ZN => n7857);
   U5395 : XNOR2_X1 port map( A => n8110, B => n7857, ZN => I2_dtemp_26_port);
   U5396 : MUX2_X1 port map( A => n8372, B => SIG_in_4_port, S => 
                           SIG_in_27_port, Z => n7862);
   U5397 : NAND2_X1 port map( A1 => n7862, A2 => SIG_in_3_port, ZN => n8055);
   U5398 : MUX2_X1 port map( A => n8373, B => n8341, S => SIG_in_27_port, Z => 
                           n8054);
   U5399 : NOR2_X1 port map( A1 => n8055, A2 => n8054, ZN => n8063);
   U5400 : MUX2_X1 port map( A => n8341, B => n2608, S => n8089, Z => n8061);
   U5401 : MUX2_X1 port map( A => n2608, B => n8365, S => n8089, Z => n8064);
   U5402 : NOR2_X1 port map( A1 => n8061, A2 => n8064, ZN => n7858);
   U5403 : NAND2_X1 port map( A1 => n8063, A2 => n7858, ZN => n8066);
   U5404 : MUX2_X1 port map( A => n8365, B => n2606, S => n8089, Z => n7867);
   U5405 : NAND2_X1 port map( A1 => n8279, A2 => n2604, ZN => n8093);
   U5406 : NOR2_X1 port map( A1 => n2606, A2 => n2605, ZN => n7859);
   U5407 : MUX2_X1 port map( A => n8371, B => SIG_in_11_port, S => n8089, Z => 
                           n8107);
   U5408 : NAND2_X1 port map( A1 => n8109, A2 => n8107, ZN => n7870);
   U5409 : MUX2_X1 port map( A => n8374, B => n2602, S => n8089, Z => n7869);
   U5410 : MUX2_X1 port map( A => n2602, B => n2601, S => n8089, Z => n8141);
   U5411 : NOR2_X1 port map( A1 => n8143, A2 => n8141, ZN => n7875);
   U5412 : MUX2_X1 port map( A => n8345, B => n8387, S => n8089, Z => n7874);
   U5413 : NAND2_X1 port map( A1 => n7875, A2 => n7874, ZN => n7873);
   U5414 : MUX2_X1 port map( A => n2600, B => n2599, S => n8089, Z => n8160);
   U5415 : NOR2_X1 port map( A1 => n7873, A2 => n8160, ZN => n7879);
   U5416 : MUX2_X1 port map( A => n8346, B => n8388, S => n8089, Z => n7878);
   U5417 : NAND2_X1 port map( A1 => n7879, A2 => n7878, ZN => n7877);
   U5418 : MUX2_X1 port map( A => n2598, B => n2597, S => n8089, Z => n8178);
   U5419 : OR2_X1 port map( A1 => n7877, A2 => n8178, ZN => n7882);
   U5420 : MUX2_X1 port map( A => n2597, B => n2596, S => n8089, Z => n7881);
   U5422 : MUX2_X1 port map( A => n2596, B => n2595, S => n8279, Z => n8199);
   U5423 : NOR2_X1 port map( A1 => n8201, A2 => n8199, ZN => n7886);
   U5424 : MUX2_X1 port map( A => n8391, B => n8348, S => n8279, Z => n7885);
   U5425 : NAND2_X1 port map( A1 => n7886, A2 => n7885, ZN => n7884);
   U5426 : MUX2_X1 port map( A => n2594, B => n2593, S => n8279, Z => n8202);
   U5427 : OR2_X1 port map( A1 => n7884, A2 => n8202, ZN => n7889);
   U5428 : MUX2_X1 port map( A => n2593, B => n2592, S => n8279, Z => n7888);
   U5430 : MUX2_X1 port map( A => n2592, B => n2591, S => n8279, Z => n8226);
   U5431 : NOR2_X1 port map( A1 => n8228, A2 => n8226, ZN => n7892);
   U5432 : MUX2_X1 port map( A => n8347, B => n8389, S => n8279, Z => n7891);
   U5433 : NAND2_X1 port map( A1 => n7892, A2 => n7891, ZN => n8261);
   U5434 : MUX2_X1 port map( A => n2590, B => n2589, S => n8279, Z => n8260);
   U5435 : NAND2_X1 port map( A1 => n8259, A2 => n8380, ZN => n8404);
   U5436 : NOR2_X1 port map( A1 => n8404, A2 => n8375, ZN => I3_SIG_out_27_port
                           );
   U5437 : AND2_X1 port map( A1 => n7861, A2 => n8354, ZN => intadd_33_A_0_port
                           );
   U5438 : OAI21_X1 port map( B1 => SIG_in_3_port, B2 => n7862, A => n8055, ZN 
                           => n7863);
   U5439 : INV_X1 port map( A => n7863, ZN => I3_SIG_out_3_port);
   U5440 : NAND2_X1 port map( A1 => n8386, A2 => n8279, ZN => n8276);
   U5441 : NOR2_X1 port map( A1 => n8276, A2 => n2577, ZN => n8278);
   U5442 : NAND2_X1 port map( A1 => n8278, A2 => EXP_in_2_port, ZN => n8275);
   U5443 : OR3_X1 port map( A1 => n8275, A2 => n8343, A3 => n8378, ZN => n8274)
                           ;
   U5444 : NOR2_X1 port map( A1 => n8274, A2 => n8384, ZN => n7864);
   U5445 : NAND2_X1 port map( A1 => n7864, A2 => n8376, ZN => n8273);
   U5446 : OR2_X1 port map( A1 => n7864, A2 => n8376, ZN => n7865);
   U5447 : AND2_X1 port map( A1 => n8273, A2 => n7865, ZN => I3_EXP_out_6_port)
                           ;
   U5448 : AND2_X1 port map( A1 => A_EXP_7_port, A2 => B_EXP_7_port, ZN => 
                           I2_EXP_pos_int);
   U5449 : OAI21_X1 port map( B1 => n8275, B2 => n8343, A => n8378, ZN => n7866
                           );
   U5450 : AND2_X1 port map( A1 => n7866, A2 => n8274, ZN => I3_EXP_out_4_port)
                           ;
   U5451 : NAND2_X1 port map( A1 => n8066, A2 => n7867, ZN => n7868);
   U5452 : AND2_X1 port map( A1 => n8092, A2 => n7868, ZN => I3_SIG_out_7_port)
                           ;
   U5453 : NAND2_X1 port map( A1 => n7870, A2 => n7869, ZN => n7871);
   U5454 : AND2_X1 port map( A1 => n8143, A2 => n7871, ZN => I3_SIG_out_11_port
                           );
   U5455 : OR2_X1 port map( A1 => n8278, A2 => EXP_in_2_port, ZN => n7872);
   U5456 : AND2_X1 port map( A1 => n8275, A2 => n7872, ZN => I3_EXP_out_2_port)
                           ;
   U5457 : OR2_X1 port map( A1 => n7875, A2 => n7874, ZN => n7876);
   U5458 : AND2_X1 port map( A1 => n7873, A2 => n7876, ZN => I3_SIG_out_13_port
                           );
   U5459 : OR2_X1 port map( A1 => n7879, A2 => n7878, ZN => n7880);
   U5460 : AND2_X1 port map( A1 => n7877, A2 => n7880, ZN => I3_SIG_out_15_port
                           );
   U5461 : NAND2_X1 port map( A1 => n7882, A2 => n7881, ZN => n7883);
   U5462 : AND2_X1 port map( A1 => n8201, A2 => n7883, ZN => I3_SIG_out_17_port
                           );
   U5463 : OR2_X1 port map( A1 => n7886, A2 => n7885, ZN => n7887);
   U5464 : AND2_X1 port map( A1 => n7884, A2 => n7887, ZN => I3_SIG_out_19_port
                           );
   U5465 : NAND2_X1 port map( A1 => n7889, A2 => n7888, ZN => n7890);
   U5466 : AND2_X1 port map( A1 => n8228, A2 => n7890, ZN => I3_SIG_out_21_port
                           );
   U5467 : OR2_X1 port map( A1 => n7892, A2 => n7891, ZN => n7893);
   U5468 : AND2_X1 port map( A1 => n8261, A2 => n7893, ZN => I3_SIG_out_23_port
                           );
   U5469 : NOR2_X1 port map( A1 => n2584, A2 => n2582, ZN => n8299);
   U5470 : NAND2_X1 port map( A1 => n8299, A2 => EXP_out_round_1_port, ZN => 
                           n8302);
   U5471 : OR2_X1 port map( A1 => n8302, A2 => n8390, ZN => n8308);
   U5472 : NAND2_X1 port map( A1 => EXP_out_round_3_port, A2 => 
                           EXP_out_round_4_port, ZN => n7894);
   U5473 : NOR2_X1 port map( A1 => n8308, A2 => n7894, ZN => n8310);
   U5474 : NAND2_X1 port map( A1 => n8310, A2 => EXP_out_round_5_port, ZN => 
                           n7913);
   U5475 : OR2_X1 port map( A1 => n7913, A2 => n2579, ZN => n7915);
   U5476 : XNOR2_X1 port map( A => n7915, B => EXP_out_round_7_port, ZN => 
                           n7917);
   U5477 : AND2_X1 port map( A1 => EXP_out_round_5_port, A2 => n8383, ZN => 
                           n7895);
   U5478 : INV_X1 port map( A => n8299, ZN => n8297);
   U5479 : NAND2_X1 port map( A1 => n2584, A2 => n2582, ZN => n8296);
   U5480 : NAND4_X1 port map( A1 => n7895, A2 => EXP_out_round_3_port, A3 => 
                           n8297, A4 => n8296, ZN => n7897);
   U5481 : NAND4_X1 port map( A1 => EXP_out_round_7_port, A2 => 
                           EXP_out_round_2_port, A3 => EXP_out_round_1_port, A4
                           => EXP_out_round_4_port, ZN => n7896);
   U5482 : OAI22_X1 port map( A1 => n7917, A2 => n2613, B1 => n7897, B2 => 
                           n7896, ZN => n8292);
   U5483 : NAND4_X1 port map( A1 => n2566, A2 => n2576, A3 => n2555, A4 => 
                           n2563, ZN => n7899);
   U5484 : NAND4_X1 port map( A1 => n2575, A2 => n2564, A3 => n2573, A4 => 
                           n2562, ZN => n7898);
   U5485 : NOR2_X1 port map( A1 => n7899, A2 => n7898, ZN => n7903);
   U5486 : NAND4_X1 port map( A1 => n2574, A2 => n2560, A3 => n2572, A4 => 
                           n2561, ZN => n7901);
   U5487 : NAND4_X1 port map( A1 => n2570, A2 => n2559, A3 => n2571, A4 => 
                           n2557, ZN => n7900);
   U5488 : NOR2_X1 port map( A1 => n7901, A2 => n7900, ZN => n7902);
   U5489 : NAND2_X1 port map( A1 => n7903, A2 => n7902, ZN => n7908);
   U5490 : AND4_X1 port map( A1 => n2569, A2 => n2558, A3 => n2556, A4 => n2568
                           , ZN => n7906);
   U5491 : NAND2_X1 port map( A1 => n2587, A2 => n2582, ZN => n7904);
   U5492 : NOR2_X1 port map( A1 => SIG_out_round_26_port, A2 => n7904, ZN => 
                           n7905);
   U5493 : NAND4_X1 port map( A1 => n7906, A2 => n7905, A3 => n2565, A4 => 
                           n8342, ZN => n7907);
   U5494 : OAI21_X1 port map( B1 => n7908, B2 => n7907, A => n2611, ZN => n7909
                           );
   U5495 : AOI21_X1 port map( B1 => n7917, B2 => EXP_neg, A => n7909, ZN => 
                           n8313);
   U5496 : OAI21_X1 port map( B1 => n8292, B2 => isINF_tab, A => n8313, ZN => 
                           n7910);
   U5497 : NAND2_X1 port map( A1 => n7910, A2 => n2567, ZN => n8315);
   U5498 : XNOR2_X1 port map( A => n8310, B => n8379, ZN => n7911);
   U5499 : AND2_X1 port map( A1 => n8313, A2 => n7911, ZN => n7912);
   U5500 : OR2_X1 port map( A1 => n8315, A2 => n7912, ZN => I4_FP_28_port);
   U5501 : NAND2_X1 port map( A1 => n7913, A2 => n2579, ZN => n7914);
   U5502 : AND3_X1 port map( A1 => n8313, A2 => n7915, A3 => n7914, ZN => n7916
                           );
   U5503 : OR2_X1 port map( A1 => n8315, A2 => n7916, ZN => I4_FP_29_port);
   U5504 : AND2_X1 port map( A1 => n8313, A2 => n7917, ZN => n7918);
   U5505 : OR2_X1 port map( A1 => n8315, A2 => n7918, ZN => I4_FP_30_port);
   U5506 : INV_X1 port map( A => n8026, ZN => n7928);
   U5507 : OAI21_X1 port map( B1 => n7920, B2 => n7928, A => n7919, ZN => n7921
                           );
   U5508 : INV_X1 port map( A => n7921, ZN => n7932);
   U5509 : INV_X1 port map( A => n7923, ZN => n8029);
   U5510 : OAI21_X1 port map( B1 => n7924, B2 => n7928, A => n8029, ZN => n7925
                           );
   U5511 : INV_X1 port map( A => n7925, ZN => n7931);
   U5512 : INV_X1 port map( A => n8032, ZN => n7926);
   U5513 : NOR2_X1 port map( A1 => n7926, A2 => n4402, ZN => n7937);
   U5514 : OR3_X1 port map( A1 => n7928, A2 => n4468, A3 => n8461, ZN => n7930)
                           ;
   U5515 : NAND4_X1 port map( A1 => n7932, A2 => n7931, A3 => n7937, A4 => 
                           n7930, ZN => n7942);
   U5516 : NAND2_X1 port map( A1 => n7934, A2 => n7933, ZN => n8028);
   U5517 : NAND2_X1 port map( A1 => n4463, A2 => n7935, ZN => n7936);
   U5518 : AOI22_X1 port map( A1 => n7937, A2 => n8028, B1 => n8032, B2 => 
                           n7936, ZN => n7941);
   U5519 : NAND2_X1 port map( A1 => n7942, A2 => n7941, ZN => n7939);
   U5520 : INV_X1 port map( A => n8428, ZN => n7938);
   U5521 : NAND2_X1 port map( A1 => n7939, A2 => n7938, ZN => n8045);
   U5522 : NAND3_X1 port map( A1 => n7942, A2 => n7941, A3 => n8428, ZN => 
                           n8044);
   U5523 : NAND2_X1 port map( A1 => n8045, A2 => n8044, ZN => n7944);
   U5524 : XNOR2_X1 port map( A => n7944, B => n7943, ZN => n8414);
   U5525 : MUX2_X1 port map( A => n7947, B => n7946, S => n7945, Z => n7948);
   U5526 : OAI21_X1 port map( B1 => n7949, B2 => n8333, A => n7948, ZN => 
                           intadd_33_B_0_port);
   U5527 : INV_X1 port map( A => n7951, ZN => n7953);
   U5528 : XNOR2_X1 port map( A => n7953, B => n7952, ZN => n7962);
   U5530 : OR2_X1 port map( A1 => n7959, A2 => n8619, ZN => n7966);
   U5531 : INV_X1 port map( A => n7959, ZN => n7955);
   U5532 : NAND3_X1 port map( A1 => n7956, A2 => n7960, A3 => n7955, ZN => 
                           n7958);
   U5533 : NAND2_X1 port map( A1 => n7962, A2 => n7959, ZN => n7957);
   U5534 : OAI211_X1 port map( C1 => n7959, C2 => n7962, A => n7958, B => n7957
                           , ZN => n7965);
   U5537 : INV_X1 port map( A => n7967, ZN => n7969);
   U5538 : NOR2_X1 port map( A1 => n7969, A2 => n7968, ZN => n7974);
   U5539 : INV_X1 port map( A => n7974, ZN => n7975);
   U5540 : NAND2_X1 port map( A1 => n7970, A2 => n7975, ZN => n7981);
   U5541 : OAI21_X1 port map( B1 => n7974, B2 => n7985, A => n7973, ZN => n7978
                           );
   U5542 : OAI21_X1 port map( B1 => n7976, B2 => n7975, A => n7984, ZN => n7977
                           );
   U5543 : NAND2_X1 port map( A1 => n7978, A2 => n7977, ZN => n7979);
   U5544 : OAI211_X1 port map( C1 => n7982, C2 => n7981, A => n7980, B => n7979
                           , ZN => n8412);
   U5545 : BUF_X1 port map( A => n7983, Z => n7995);
   U5546 : XNOR2_X1 port map( A => n7985, B => n7984, ZN => n7994);
   U5547 : NAND2_X1 port map( A1 => n7986, A2 => n4459, ZN => n7987);
   U5549 : INV_X1 port map( A => n8563, ZN => n7991);
   U5551 : NAND2_X1 port map( A1 => n7991, A2 => n8614, ZN => n7992);
   U5553 : INV_X1 port map( A => n8280, ZN => n7996);
   U5554 : NAND2_X1 port map( A1 => n7997, A2 => n7996, ZN => n8001);
   U5555 : INV_X1 port map( A => I1_I1_N13, ZN => n7998);
   U5556 : NAND2_X1 port map( A1 => n7999, A2 => n7998, ZN => n8000);
   U5557 : AOI21_X1 port map( B1 => n8001, B2 => n8000, A => n8284, ZN => 
                           I1_isZ_tab_int);
   U5558 : XNOR2_X1 port map( A => n381, B => n8002, ZN => n8006);
   U5559 : MUX2_X1 port map( A => n8459, B => n8434, S => n8393, Z => n8005);
   U5560 : OAI21_X1 port map( B1 => n8007, B2 => n8006, A => n8005, ZN => 
                           intadd_33_CI);
   U5561 : OAI21_X1 port map( B1 => n8010, B2 => n8009, A => n8008, ZN => n8011
                           );
   U5562 : INV_X1 port map( A => n8011, ZN => intadd_33_A_1_port);
   U5563 : MUX2_X1 port map( A => n4975, B => n8012, S => n8401, Z => n8013);
   U5564 : INV_X1 port map( A => n8013, ZN => n8015);
   U5565 : MUX2_X1 port map( A => n5878, B => n6102, S => n8350, Z => n8014);
   U5566 : NAND2_X1 port map( A1 => n8015, A2 => n8014, ZN => 
                           intadd_33_B_1_port);
   U5567 : XNOR2_X1 port map( A => n8017, B => n8016, ZN => n8019);
   U5568 : XNOR2_X1 port map( A => n8018, B => n8019, ZN => n8408);
   U5569 : NAND2_X1 port map( A1 => n8021, A2 => n8020, ZN => n8024);
   U5570 : INV_X1 port map( A => n8022, ZN => n8023);
   U5571 : XNOR2_X1 port map( A => n8024, B => n8023, ZN => intadd_33_B_2_port)
                           ;
   U5573 : NAND2_X1 port map( A1 => n8027, A2 => n8026, ZN => n8030);
   U5574 : AOI21_X1 port map( B1 => n8030, B2 => n8029, A => n8028, ZN => n8039
                           );
   U5575 : OAI21_X1 port map( B1 => n8039, B2 => n4402, A => n7935, ZN => n8035
                           );
   U5576 : AND2_X1 port map( A1 => n4463, A2 => n8032, ZN => n8034);
   U5577 : XNOR2_X1 port map( A => n8035, B => n8034, ZN => I2_dtemp_23_port);
   U5578 : XNOR2_X1 port map( A => n8037, B => n8036, ZN => n8038);
   U5579 : XNOR2_X1 port map( A => n8039, B => n8038, ZN => n8407);
   U5580 : INV_X1 port map( A => n8040, ZN => n8041);
   U5581 : NAND2_X1 port map( A1 => n8044, A2 => n8041, ZN => n8047);
   U5582 : INV_X1 port map( A => n8042, ZN => n8043);
   U5583 : NAND2_X1 port map( A1 => n8044, A2 => n8043, ZN => n8046);
   U5584 : NAND3_X1 port map( A1 => n8047, A2 => n8046, A3 => n8045, ZN => 
                           n8053);
   U5585 : OAI21_X1 port map( B1 => n8050, B2 => n8449, A => n8048, ZN => n8051
                           );
   U5586 : INV_X1 port map( A => n8051, ZN => n8052);
   U5587 : XNOR2_X1 port map( A => n8053, B => n8052, ZN => n8413);
   U5588 : AND2_X1 port map( A1 => n8055, A2 => n8054, ZN => n8056);
   U5589 : NOR2_X1 port map( A1 => n8063, A2 => n8056, ZN => I3_SIG_out_4_port)
                           ;
   U5590 : XNOR2_X1 port map( A => n8061, B => n8063, ZN => I3_SIG_out_5_port);
   U5591 : NAND2_X1 port map( A1 => n8444, A2 => n8490, ZN => n8060);
   U5592 : INV_X1 port map( A => n8079, ZN => n8058);
   U5593 : NAND2_X1 port map( A1 => n8058, A2 => n8075, ZN => n8059);
   U5594 : XNOR2_X1 port map( A => n8060, B => n8059, ZN => I2_dtemp_27_port);
   U5595 : INV_X1 port map( A => n8061, ZN => n8062);
   U5596 : NAND2_X1 port map( A1 => n8063, A2 => n8062, ZN => n8065);
   U5597 : NAND2_X1 port map( A1 => n8065, A2 => n8064, ZN => n8067);
   U5598 : AND2_X1 port map( A1 => n8067, A2 => n8066, ZN => I3_SIG_out_6_port)
                           ;
   U5599 : XNOR2_X1 port map( A => n4444, B => n8077, ZN => n8072);
   U5600 : OAI21_X1 port map( B1 => n8079, B2 => n8490, A => n8075, ZN => n8068
                           );
   U5601 : INV_X1 port map( A => n8068, ZN => n8069);
   U5602 : OAI21_X1 port map( B1 => n8444, B2 => n8079, A => n8069, ZN => n8071
                           );
   U5603 : NAND2_X1 port map( A1 => n8071, A2 => n8072, ZN => n8070);
   U5604 : OAI21_X1 port map( B1 => n8072, B2 => n8071, A => n8070, ZN => 
                           I2_dtemp_28_port);
   U5605 : NAND2_X1 port map( A1 => n8444, A2 => n4533, ZN => n8084);
   U5606 : INV_X1 port map( A => n4444, ZN => n8081);
   U5607 : INV_X1 port map( A => n8077, ZN => n8078);
   U5608 : OAI21_X1 port map( B1 => n8079, B2 => n8081, A => n8078, ZN => n8080
                           );
   U5609 : NAND2_X1 port map( A1 => n8084, A2 => n8083, ZN => n8088);
   U5610 : XNOR2_X1 port map( A => n8594, B => n8085, ZN => n8087);
   U5611 : XNOR2_X1 port map( A => n8088, B => n8087, ZN => n8406);
   U5612 : MUX2_X1 port map( A => n2606, B => n2605, S => n8089, Z => n8091);
   U5613 : INV_X1 port map( A => n8091, ZN => n8090);
   U5614 : XNOR2_X1 port map( A => n8092, B => n8090, ZN => I3_SIG_out_8_port);
   U5615 : NOR2_X1 port map( A1 => n8092, A2 => n8091, ZN => n8095);
   U5616 : OAI21_X1 port map( B1 => n8279, B2 => n8381, A => n8093, ZN => n8094
                           );
   U5617 : XNOR2_X1 port map( A => n8095, B => n8094, ZN => I3_SIG_out_9_port);
   U5618 : NOR2_X1 port map( A1 => n8096, A2 => n4399, ZN => n8122);
   U5619 : NAND2_X1 port map( A1 => n8444, A2 => n8122, ZN => n8102);
   U5620 : AOI22_X1 port map( A1 => n8100, A2 => n8099, B1 => n8098, B2 => 
                           n8584, ZN => n8101);
   U5621 : NAND2_X1 port map( A1 => n8102, A2 => n8101, ZN => n8106);
   U5622 : AND2_X1 port map( A1 => n8104, A2 => n8123, ZN => n8105);
   U5623 : XNOR2_X1 port map( A => n8106, B => n8105, ZN => I2_dtemp_31_port);
   U5624 : INV_X1 port map( A => n8107, ZN => n8108);
   U5625 : XNOR2_X1 port map( A => n8109, B => n8108, ZN => I3_SIG_out_10_port)
                           ;
   U5626 : NAND3_X1 port map( A1 => n8110, A2 => n8122, A3 => n8104, ZN => 
                           n8114);
   U5627 : INV_X1 port map( A => n8104, ZN => n8137);
   U5628 : NOR2_X1 port map( A1 => n4399, A2 => n8137, ZN => n8112);
   U5629 : AOI21_X1 port map( B1 => n4459, B2 => n8112, A => n8111, ZN => n8113
                           );
   U5630 : NAND2_X1 port map( A1 => n8114, A2 => n8113, ZN => n8119);
   U5632 : XOR2_X1 port map( A => n8450, B => n8117, Z => n8118);
   U5633 : XNOR2_X1 port map( A => n8119, B => n8118, ZN => n8405);
   U5634 : INV_X1 port map( A => n4459, ZN => n8125);
   U5635 : NAND2_X1 port map( A1 => n8121, A2 => n8122, ZN => n8124);
   U5636 : AND2_X1 port map( A1 => n8126, A2 => n4485, ZN => n8130);
   U5637 : INV_X1 port map( A => n8130, ZN => n8132);
   U5638 : AND2_X1 port map( A1 => n8132, A2 => n4426, ZN => n8136);
   U5639 : INV_X1 port map( A => n8136, ZN => n8140);
   U5640 : NAND2_X1 port map( A1 => n8130, A2 => n4426, ZN => n8135);
   U5642 : NAND2_X1 port map( A1 => n8466, A2 => n8132, ZN => n8134);
   U5643 : AOI22_X1 port map( A1 => n8137, A2 => n8136, B1 => n8135, B2 => 
                           n8134, ZN => n8138);
   U5644 : OAI211_X1 port map( C1 => n4503, C2 => n8140, A => n8139, B => n8138
                           , ZN => I2_dtemp_33_port);
   U5645 : INV_X1 port map( A => n8141, ZN => n8142);
   U5646 : XNOR2_X1 port map( A => n8143, B => n8142, ZN => I3_SIG_out_12_port)
                           ;
   U5647 : NOR2_X1 port map( A1 => n7727, A2 => n8147, ZN => n8148);
   U5648 : OR2_X1 port map( A1 => n4428, A2 => n8148, ZN => n8154);
   U5649 : INV_X1 port map( A => n8162, ZN => n8155);
   U5650 : NAND2_X1 port map( A1 => n8155, A2 => n4498, ZN => n8150);
   U5652 : NAND3_X1 port map( A1 => n8154, A2 => n4498, A3 => n4485, ZN => 
                           n8156);
   U5653 : OAI21_X1 port map( B1 => n8174, B2 => n8156, A => n8155, ZN => n8159
                           );
   U5654 : AND2_X1 port map( A1 => n7597, A2 => n8580, ZN => n8158);
   U5655 : XNOR2_X1 port map( A => n8159, B => n8158, ZN => n8410);
   U5656 : INV_X1 port map( A => n8160, ZN => n8161);
   U5657 : XNOR2_X1 port map( A => n7873, B => n8161, ZN => I3_SIG_out_14_port)
                           ;
   U5658 : NAND2_X1 port map( A1 => n8192, A2 => n4500, ZN => n8164);
   U5659 : NAND2_X1 port map( A1 => n8162, A2 => n8580, ZN => n8163);
   U5660 : AND2_X1 port map( A1 => n7597, A2 => n8163, ZN => n8170);
   U5661 : OAI21_X1 port map( B1 => n8174, B2 => n8164, A => n8170, ZN => n8166
                           );
   U5662 : XNOR2_X1 port map( A => n8166, B => n8165, ZN => n8409);
   U5663 : INV_X1 port map( A => n7606, ZN => n8167);
   U5664 : NAND3_X1 port map( A1 => n8192, A2 => n4500, A3 => n8167, ZN => 
                           n8173);
   U5665 : INV_X1 port map( A => n8168, ZN => n8169);
   U5666 : OAI21_X1 port map( B1 => n8170, B2 => n7606, A => n8169, ZN => n8171
                           );
   U5667 : INV_X1 port map( A => n8171, ZN => n8172);
   U5668 : OAI21_X1 port map( B1 => n8174, B2 => n8173, A => n8172, ZN => n8177
                           );
   U5669 : AND2_X1 port map( A1 => n8175, A2 => n7377, ZN => n8176);
   U5670 : XNOR2_X1 port map( A => n8177, B => n8176, ZN => I2_dtemp_37_port);
   U5671 : INV_X1 port map( A => n8178, ZN => n8179);
   U5672 : XNOR2_X1 port map( A => n7877, B => n8179, ZN => I3_SIG_out_16_port)
                           ;
   U5673 : INV_X1 port map( A => n8186, ZN => n8182);
   U5674 : XNOR2_X1 port map( A => n8181, B => n8180, ZN => n8185);
   U5675 : NAND2_X1 port map( A1 => n8182, A2 => n8185, ZN => n8198);
   U5676 : NOR2_X1 port map( A1 => n8189, A2 => n8185, ZN => n8183);
   U5677 : NAND4_X1 port map( A1 => n8184, A2 => n8192, A3 => n8183, A4 => 
                           n8480, ZN => n8196);
   U5678 : NOR2_X1 port map( A1 => n8184, A2 => n8198, ZN => n8194);
   U5679 : INV_X1 port map( A => n8185, ZN => n8187);
   U5680 : AND2_X1 port map( A1 => n8186, A2 => n8187, ZN => n8190);
   U5681 : NAND2_X1 port map( A1 => n8189, A2 => n8187, ZN => n8188);
   U5682 : OAI21_X1 port map( B1 => n8190, B2 => n8189, A => n8188, ZN => n8191
                           );
   U5683 : OAI21_X1 port map( B1 => n8192, B2 => n8198, A => n8191, ZN => n8193
                           );
   U5684 : NOR2_X1 port map( A1 => n8194, A2 => n8193, ZN => n8195);
   U5685 : OAI211_X1 port map( C1 => n8198, C2 => n8480, A => n8195, B => n8196
                           , ZN => I2_dtemp_38_port);
   U5686 : INV_X1 port map( A => n8199, ZN => n8200);
   U5687 : XNOR2_X1 port map( A => n8201, B => n8200, ZN => I3_SIG_out_18_port)
                           ;
   U5688 : INV_X1 port map( A => n8202, ZN => n8203);
   U5689 : XNOR2_X1 port map( A => n7884, B => n8203, ZN => I3_SIG_out_20_port)
                           ;
   U5691 : NAND2_X1 port map( A1 => n8206, A2 => n8205, ZN => n8216);
   U5692 : NAND3_X1 port map( A1 => n8208, A2 => n8207, A3 => n8216, ZN => 
                           n8239);
   U5694 : NAND2_X1 port map( A1 => n8252, A2 => n8601, ZN => n8237);
   U5695 : OR2_X1 port map( A1 => n8239, A2 => n4399, ZN => n8211);
   U5696 : NOR2_X1 port map( A1 => n8212, A2 => n8211, ZN => n8254);
   U5697 : NAND2_X1 port map( A1 => n8254, A2 => n4459, ZN => n8235);
   U5698 : INV_X1 port map( A => n8240, ZN => n8243);
   U5699 : XNOR2_X1 port map( A => n7711, B => n8243, ZN => n8223);
   U5700 : INV_X1 port map( A => n8223, ZN => n8220);
   U5701 : INV_X1 port map( A => n8213, ZN => n8217);
   U5702 : INV_X1 port map( A => n8214, ZN => n8215);
   U5703 : AOI21_X1 port map( B1 => n8217, B2 => n8216, A => n8215, ZN => n8248
                           );
   U5704 : NAND2_X1 port map( A1 => n8229, A2 => n8248, ZN => n8219);
   U5705 : NAND2_X1 port map( A1 => n8239, A2 => n8248, ZN => n8218);
   U5706 : NAND2_X1 port map( A1 => n8219, A2 => n8218, ZN => n8221);
   U5707 : NAND4_X1 port map( A1 => n8237, A2 => n8235, A3 => n8220, A4 => 
                           n8221, ZN => n8225);
   U5708 : INV_X1 port map( A => n8221, ZN => n8222);
   U5709 : NAND2_X1 port map( A1 => n8222, A2 => n8223, ZN => n8224);
   U5710 : INV_X1 port map( A => n8226, ZN => n8227);
   U5711 : XNOR2_X1 port map( A => n8228, B => n8227, ZN => I3_SIG_out_22_port)
                           ;
   U5712 : INV_X1 port map( A => n8229, ZN => n8251);
   U5713 : INV_X1 port map( A => n8239, ZN => n8234);
   U5714 : NAND2_X1 port map( A1 => n8231, A2 => n8230, ZN => n8241);
   U5715 : NAND3_X1 port map( A1 => n8248, A2 => n8232, A3 => n8241, ZN => 
                           n8233);
   U5716 : AOI21_X1 port map( B1 => n8251, B2 => n8234, A => n8233, ZN => n8236
                           );
   U5717 : NAND3_X1 port map( A1 => n8237, A2 => n8236, A3 => n8235, ZN => 
                           n8258);
   U5718 : INV_X1 port map( A => n8241, ZN => n8244);
   U5719 : AND2_X1 port map( A1 => n8238, A2 => n8244, ZN => n8253);
   U5720 : INV_X1 port map( A => n8253, ZN => n8247);
   U5721 : NOR2_X1 port map( A1 => n8239, A2 => n8247, ZN => n8250);
   U5722 : NAND2_X1 port map( A1 => n8241, A2 => n8240, ZN => n8242);
   U5723 : AND2_X1 port map( A1 => n8242, A2 => n7711, ZN => n8246);
   U5724 : AOI21_X1 port map( B1 => n8244, B2 => n8243, A => n7711, ZN => n8245
                           );
   U5725 : OAI22_X1 port map( A1 => n8248, A2 => n8247, B1 => n8246, B2 => 
                           n8245, ZN => n8249);
   U5726 : AOI21_X1 port map( B1 => n8251, B2 => n8250, A => n8249, ZN => n8257
                           );
   U5727 : NAND3_X1 port map( A1 => n8252, A2 => n8601, A3 => n8253, ZN => 
                           n8256);
   U5728 : NAND3_X1 port map( A1 => n4459, A2 => n8254, A3 => n8253, ZN => 
                           n8255);
   U5729 : NAND4_X1 port map( A1 => n8258, A2 => n8257, A3 => n8256, A4 => 
                           n8255, ZN => I2_dtemp_44_port);
   U5730 : AND2_X1 port map( A1 => n8261, A2 => n8260, ZN => n8262);
   U5731 : NOR2_X1 port map( A1 => n8259, A2 => n8262, ZN => I3_SIG_out_24_port
                           );
   U5732 : MUX2_X1 port map( A => n2589, B => n8375, S => n8279, Z => n8263);
   U5733 : XNOR2_X1 port map( A => n8259, B => n8263, ZN => I3_SIG_out_25_port)
                           ;
   U5734 : NAND4_X1 port map( A1 => A_EXP_2_port, A2 => A_EXP_3_port, A3 => 
                           A_EXP_4_port, A4 => A_EXP_5_port, ZN => n8266);
   U5735 : NAND3_X1 port map( A1 => A_EXP_6_port, A2 => A_EXP_0_port, A3 => 
                           A_EXP_1_port, ZN => n8265);
   U5736 : NOR2_X1 port map( A1 => A_EXP_7_port, A2 => B_EXP_7_port, ZN => 
                           n8264);
   U5737 : OAI21_X1 port map( B1 => n8266, B2 => n8265, A => n8264, ZN => n8270
                           );
   U5738 : NAND4_X1 port map( A1 => B_EXP_1_port, A2 => B_EXP_2_port, A3 => 
                           B_EXP_4_port, A4 => B_EXP_5_port, ZN => n8268);
   U5739 : NAND3_X1 port map( A1 => B_EXP_0_port, A2 => B_EXP_6_port, A3 => 
                           B_EXP_3_port, ZN => n8267);
   U5740 : NOR2_X1 port map( A1 => n8268, A2 => n8267, ZN => n8269);
   U5741 : NOR2_X1 port map( A1 => n8270, A2 => n8269, ZN => I2_N0);
   U5742 : NAND2_X1 port map( A1 => n8382, A2 => n8344, ZN => intadd_2_CI);
   U5743 : XOR2_X1 port map( A => A_EXP_7_port, B => B_EXP_7_port, Z => n8271);
   U5744 : XNOR2_X1 port map( A => intadd_2_n1, B => n8271, ZN => n374);
   U5745 : NAND2_X1 port map( A1 => B_EXP_0_port, A2 => A_EXP_0_port, ZN => 
                           n8272);
   U5746 : NAND2_X1 port map( A1 => intadd_2_CI, A2 => n8272, ZN => 
                           I2_mw_I4sum_0_port);
   U5747 : XNOR2_X1 port map( A => n8273, B => EXP_in_7_port, ZN => 
                           I3_EXP_out_7_port);
   U5748 : XNOR2_X1 port map( A => n8274, B => EXP_in_5_port, ZN => 
                           I3_EXP_out_5_port);
   U5749 : XNOR2_X1 port map( A => n8275, B => EXP_in_3_port, ZN => 
                           I3_EXP_out_3_port);
   U5750 : AND2_X1 port map( A1 => n8276, A2 => n2577, ZN => n8277);
   U5751 : NOR2_X1 port map( A1 => n8278, A2 => n8277, ZN => I3_EXP_out_1_port)
                           ;
   U5752 : XNOR2_X1 port map( A => n8279, B => n2583, ZN => I3_EXP_out_0_port);
   U5753 : NAND2_X1 port map( A1 => n8281, A2 => n8280, ZN => n8286);
   U5754 : NAND2_X1 port map( A1 => n8283, A2 => n8282, ZN => n8285);
   U5755 : MUX2_X1 port map( A => n8286, B => n8285, S => n8284, Z => n8288);
   U5756 : NAND2_X1 port map( A1 => n8288, A2 => n8287, ZN => I1_isNaN_int);
   U5757 : INV_X1 port map( A => n8313, ZN => n8289);
   U5758 : OAI22_X1 port map( A1 => n2565, A2 => n8290, B1 => n8291, B2 => 
                           n2587, ZN => I4_FP_0_port);
   U5759 : OAI22_X1 port map( A1 => n2565, A2 => n8291, B1 => n8290, B2 => 
                           n2556, ZN => I4_FP_1_port);
   U5760 : OAI22_X1 port map( A1 => n2568, A2 => n8290, B1 => n8291, B2 => 
                           n2556, ZN => I4_FP_2_port);
   U5761 : OAI22_X1 port map( A1 => n2557, A2 => n8290, B1 => n8291, B2 => 
                           n2568, ZN => I4_FP_3_port);
   U5762 : OAI22_X1 port map( A1 => n2557, A2 => n8291, B1 => n8290, B2 => 
                           n2569, ZN => I4_FP_4_port);
   U5763 : OAI22_X1 port map( A1 => n2558, A2 => n8290, B1 => n8291, B2 => 
                           n2569, ZN => I4_FP_5_port);
   U5764 : OAI22_X1 port map( A1 => n2570, A2 => n8290, B1 => n8291, B2 => 
                           n2558, ZN => I4_FP_6_port);
   U5765 : OAI22_X1 port map( A1 => n2559, A2 => n8290, B1 => n8291, B2 => 
                           n2570, ZN => I4_FP_7_port);
   U5766 : OAI22_X1 port map( A1 => n2571, A2 => n8290, B1 => n8291, B2 => 
                           n2559, ZN => I4_FP_8_port);
   U5767 : OAI22_X1 port map( A1 => n2571, A2 => n8291, B1 => n8290, B2 => 
                           n2560, ZN => I4_FP_9_port);
   U5768 : OAI22_X1 port map( A1 => n2572, A2 => n8290, B1 => n8291, B2 => 
                           n2560, ZN => I4_FP_10_port);
   U5769 : OAI22_X1 port map( A1 => n2561, A2 => n8290, B1 => n8291, B2 => 
                           n2572, ZN => I4_FP_11_port);
   U5770 : OAI22_X1 port map( A1 => n2561, A2 => n8291, B1 => n8290, B2 => 
                           n2573, ZN => I4_FP_12_port);
   U5771 : OAI22_X1 port map( A1 => n2562, A2 => n8290, B1 => n8291, B2 => 
                           n2573, ZN => I4_FP_13_port);
   U5772 : OAI22_X1 port map( A1 => n2574, A2 => n8290, B1 => n8291, B2 => 
                           n2562, ZN => I4_FP_14_port);
   U5773 : OAI22_X1 port map( A1 => n2574, A2 => n8291, B1 => n8290, B2 => 
                           n2563, ZN => I4_FP_15_port);
   U5774 : OAI22_X1 port map( A1 => n2575, A2 => n8290, B1 => n8291, B2 => 
                           n2563, ZN => I4_FP_16_port);
   U5775 : OAI22_X1 port map( A1 => n2564, A2 => n8290, B1 => n8291, B2 => 
                           n2575, ZN => I4_FP_17_port);
   U5776 : OAI22_X1 port map( A1 => n2564, A2 => n8291, B1 => n8290, B2 => 
                           n2576, ZN => I4_FP_18_port);
   U5777 : OAI22_X1 port map( A1 => n2555, A2 => n8290, B1 => n8291, B2 => 
                           n2576, ZN => I4_FP_19_port);
   U5778 : OAI22_X1 port map( A1 => n2555, A2 => n8291, B1 => n8290, B2 => 
                           n2566, ZN => I4_FP_20_port);
   U5779 : OAI22_X1 port map( A1 => n2566, A2 => n8291, B1 => n8290, B2 => 
                           n8342, ZN => I4_FP_21_port);
   U5780 : INV_X1 port map( A => n8292, ZN => n8294);
   U5781 : MUX2_X1 port map( A => SIG_out_round_26_port, B => 
                           SIG_out_round_25_port, S => n2582, Z => n8293);
   U5782 : NAND4_X1 port map( A1 => n8294, A2 => n8313, A3 => n8385, A4 => 
                           n8293, ZN => n8295);
   U5783 : NAND2_X1 port map( A1 => n8295, A2 => n2567, ZN => I4_FP_22_port);
   U5784 : AND3_X1 port map( A1 => n8313, A2 => n8297, A3 => n8296, ZN => n8298
                           );
   U5785 : OR2_X1 port map( A1 => n8315, A2 => n8298, ZN => I4_FP_23_port);
   U5786 : INV_X1 port map( A => n8315, ZN => n8301);
   U5787 : OAI211_X1 port map( C1 => n8299, C2 => EXP_out_round_1_port, A => 
                           n8313, B => n8302, ZN => n8300);
   U5788 : NAND2_X1 port map( A1 => n8301, A2 => n8300, ZN => I4_FP_24_port);
   U5789 : INV_X1 port map( A => n8302, ZN => n8303);
   U5790 : OAI211_X1 port map( C1 => EXP_out_round_2_port, C2 => n8303, A => 
                           n8313, B => n8308, ZN => n8304);
   U5791 : INV_X1 port map( A => n8304, ZN => n8305);
   U5792 : OR2_X1 port map( A1 => n8315, A2 => n8305, ZN => I4_FP_25_port);
   U5793 : XNOR2_X1 port map( A => n8308, B => EXP_out_round_3_port, ZN => 
                           n8306);
   U5794 : AND2_X1 port map( A1 => n8313, A2 => n8306, ZN => n8307);
   U5795 : OR2_X1 port map( A1 => n8315, A2 => n8307, ZN => I4_FP_26_port);
   U5796 : INV_X1 port map( A => n8308, ZN => n8309);
   U5797 : AOI21_X1 port map( B1 => n8309, B2 => EXP_out_round_3_port, A => 
                           EXP_out_round_4_port, ZN => n8311);
   U5798 : NOR2_X1 port map( A1 => n8311, A2 => n8310, ZN => n8312);
   U5799 : AND2_X1 port map( A1 => n8313, A2 => n8312, ZN => n8314);
   U5800 : OR2_X1 port map( A1 => n8315, A2 => n8314, ZN => I4_FP_27_port);
   U5801 : INV_X1 port map( A => FP_B(31), ZN => n8316);
   U5802 : XNOR2_X1 port map( A => n8316, B => FP_A(31), ZN => I1_SIGN_out_int)
                           ;
   I1_B_EXP_reg_3_inst : DFF_X1 port map( D => FP_B(26), CK => clk, Q => 
                           B_EXP_3_port, QN => n_1142);
   I2_EXP_in_reg_4_inst : DFF_X1 port map( D => n8323, CK => clk, Q => n8378, 
                           QN => n_1143);
   I2_EXP_in_tmp_reg_4_inst : DFF_X1 port map( D => I2_mw_I4sum_4_port, CK => 
                           clk, Q => n_1144, QN => n8323);
   I2_SIG_in_reg_20_inst : DFF_X1 port map( D => I2_SIG_in_int_20_port, CK => 
                           clk, Q => n8348, QN => n2594);
   I1_B_SIG_reg_2_inst : DFF_X1 port map( D => FP_B(2), CK => clk, Q => n8396, 
                           QN => n381);
   I2_SIG_in_reg_2_inst : SDFF_X1 port map( D => I2_SIG_in_int_2_port, SI => 
                           n8520, SE => n8520, CK => clk, Q => n8372, QN => 
                           n_1145);
   I2_SIG_in_reg_27_inst : SDFF_X1 port map( D => I2_SIG_in_int_27_port, SI => 
                           n8518, SE => n8518, CK => clk, Q => SIG_in_27_port, 
                           QN => n_1146);
   U5149 : BUF_X2 port map( A => n8121, Z => n8110);
   U1794 : BUF_X1 port map( A => n6420, Z => n6391);
   U1809 : AND2_X2 port map( A1 => n8154, A2 => n4485, ZN => n8192);
   U1886 : BUF_X2 port map( A => n5867, Z => n7559);
   U1749 : NAND2_X1 port map( A1 => n8208, A2 => n7732, ZN => n7728);
   U2400 : NOR2_X1 port map( A1 => n8335, A2 => n389, ZN => n6738);
   U1949 : OR2_X1 port map( A1 => n8355, A2 => n164, ZN => n5760);
   U2250 : BUF_X2 port map( A => n391, Z => n5879);
   U3196 : BUF_X1 port map( A => n7090, Z => n7696);
   U2572 : OAI211_X1 port map( C1 => n395, C2 => n8593, A => n4726, B => n4725,
                           ZN => n4954);
   U1746 : MUX2_X1 port map( A => n4487, B => n7325, S => n359, Z => n6399);
   U2367 : NAND2_X1 port map( A1 => n4550, A2 => n4549, ZN => n4554);
   U1982 : NOR2_X1 port map( A1 => n8462, A2 => n4553, ZN => n4423);
   U1795 : OR2_X1 port map( A1 => n5394, A2 => n5393, ZN => n5598);
   U1774 : AND2_X1 port map( A1 => n4354, A2 => n4353, ZN => n7039);
   U1737 : OR2_X1 port map( A1 => n7870, A2 => n7869, ZN => n8143);
   U1770 : AND2_X1 port map( A1 => n5485, A2 => n5484, ZN => n5678);
   U2906 : XNOR2_X1 port map( A => n5071, B => n5202, ZN => n5182);
   U5421 : OR2_X1 port map( A1 => n7882, A2 => n7881, ZN => n8201);
   U1733 : NAND2_X1 port map( A1 => n6340, A2 => n6339, ZN => n6548);
   U1741 : OR2_X1 port map( A1 => n4506, A2 => n5253, ZN => n5263);
   U5429 : OR2_X1 port map( A1 => n7889, A2 => n7888, ZN => n8228);
   U1816 : BUF_X1 port map( A => n8031, Z => n4402);
   U2107 : INV_X2 port map( A => n8398, ZN => n4514);
   U1895 : INV_X1 port map( A => n5302, ZN => n5303);
   U2021 : INV_X2 port map( A => n5872, ZN => n6887);
   U1857 : OR2_X1 port map( A1 => n6436, A2 => n6435, ZN => n6483);
   U2078 : AOI21_X1 port map( B1 => n6855, B2 => n6856, A => n6854, ZN => n6869
                           );
   U3870 : NOR2_X2 port map( A1 => n7619, A2 => n7620, ZN => n8209);
   U1968 : OR2_X2 port map( A1 => n6775, A2 => n6774, ZN => n6982);
   U2340 : NAND2_X2 port map( A1 => n5051, A2 => n5854, ZN => n6888);
   U2353 : NAND3_X2 port map( A1 => n5883, A2 => n5854, A3 => A_SIG_10_port, ZN
                           => n4607);
   I2_prod_tmp_reg_41_inst : DFF_X1 port map( D => I2_dtemp_41_port, CK => clk,
                           Q => I2_SIG_in_int_21_port, QN => n_1147);
   I2_prod_tmp_reg_31_inst : DFF_X1 port map( D => I2_dtemp_31_port, CK => clk,
                           Q => I2_SIG_in_int_11_port, QN => n_1148);
   U1731 : OR2_X2 port map( A1 => n6617, A2 => n6616, ZN => n6721);
   U1740 : OAI22_X1 port map( A1 => n5571, A2 => n5575, B1 => n5573, B2 => 
                           n5570, ZN => n7923);
   U1759 : MUX2_X1 port map( A => n6812, B => n8593, S => n8329, Z => n6693);
   U1761 : MUX2_X1 port map( A => n7123, B => n6812, S => n2638, Z => n4550);
   U1764 : CLKBUF_X1 port map( A => n8025, Z => n8027);
   U1769 : AND4_X2 port map( A1 => n6085, A2 => n8048, A3 => n8032, A4 => n6084
                           , ZN => n6086);
   U1771 : OAI21_X2 port map( B1 => n4512, B2 => n6882, A => n6883, ZN => n7062
                           );
   U1777 : CLKBUF_X1 port map( A => n7972, Z => n7982);
   U1813 : BUF_X1 port map( A => n8073, Z => n8490);
   U1825 : OR2_X1 port map( A1 => n8116, A2 => n8115, ZN => n8131);
   U1826 : NAND2_X1 port map( A1 => n8426, A2 => n8425, ZN => n6523);
   U1827 : OAI21_X1 port map( B1 => n8569, B2 => n6521, A => n6522, ZN => n8426
                           );
   U1837 : AOI21_X1 port map( B1 => n6601, B2 => n6949, A => n8416, ZN => n6959
                           );
   U1851 : AND2_X1 port map( A1 => n5493, A2 => n5492, ZN => n5669);
   U1855 : NOR2_X1 port map( A1 => n7034, A2 => n7035, ZN => n7038);
   U1859 : AND2_X1 port map( A1 => n8424, A2 => n8422, ZN => n5440);
   U1887 : OR2_X1 port map( A1 => n5865, A2 => n4528, ZN => n6174);
   U1891 : AND2_X1 port map( A1 => n5848, A2 => n4538, ZN => n4561);
   U1930 : INV_X1 port map( A => n8399, ZN => n8503);
   U1947 : INV_X1 port map( A => n4553, ZN => n8421);
   U1956 : NAND2_X1 port map( A1 => n4606, A2 => n4605, ZN => n4621);
   U1961 : NAND2_X1 port map( A1 => n6112, A2 => n6111, ZN => n6121);
   U1969 : AOI21_X1 port map( B1 => n7216, B2 => n8349, A => n7036, ZN => n4354
                           );
   U1977 : OAI22_X1 port map( A1 => n6851, A2 => n6850, B1 => n6849, B2 => 
                           n6848, ZN => n6867);
   U1998 : OR2_X1 port map( A1 => n4618, A2 => n4617, ZN => n4689);
   U1999 : AOI22_X1 port map( A1 => n5131, A2 => n5130, B1 => n5129, B2 => 
                           n5128, ZN => n5156);
   U2004 : XNOR2_X1 port map( A => n5292, B => n5681, ZN => n5470);
   U2009 : OR2_X1 port map( A1 => n7205, A2 => n7206, ZN => n7319);
   U2049 : NAND2_X1 port map( A1 => n8569, A2 => n6521, ZN => n8425);
   U2072 : CLKBUF_X1 port map( A => n6077, Z => n8467);
   U2100 : XNOR2_X1 port map( A => n5540, B => n5539, ZN => n5827);
   U2104 : OAI21_X1 port map( B1 => n7571, B2 => n7574, A => n7572, ZN => n7712
                           );
   U2106 : OR2_X1 port map( A1 => n4413, A2 => n6556, ZN => n6559);
   U2114 : OAI22_X1 port map( A1 => n7986, A2 => n8615, B1 => n7740, B2 => 
                           n7739, ZN => n4445);
   U2144 : CLKBUF_X1 port map( A => n8116, Z => n8117);
   U2160 : NOR2_X1 port map( A1 => n7376, A2 => n7375, ZN => n8168);
   U2183 : AOI21_X1 port map( B1 => n4447, B2 => n8209, A => n8239, ZN => n8252
                           );
   U2197 : OAI21_X1 port map( B1 => n8144, B2 => n8145, A => n8152, ZN => n8174
                           );
   U2218 : AND2_X1 port map( A1 => n6258, A2 => n6257, ZN => n8415);
   U2220 : AND2_X1 port map( A1 => n6602, A2 => n6948, ZN => n8416);
   U2225 : NAND2_X1 port map( A1 => n8420, A2 => n8417, ZN => n6417);
   U2242 : NOR2_X1 port map( A1 => n8419, A2 => n8418, ZN => n8417);
   U2251 : INV_X1 port map( A => n6411, ZN => n8418);
   U2307 : INV_X1 port map( A => n6412, ZN => n8419);
   U2308 : NAND2_X1 port map( A1 => n6413, A2 => n6409, ZN => n8420);
   U2309 : INV_X1 port map( A => n4621, ZN => n4619);
   U2310 : NAND3_X1 port map( A1 => n6984, A2 => n6982, A3 => n6983, ZN => 
                           n8116);
   U2311 : NAND2_X1 port map( A1 => n4554, A2 => n8421, ZN => n4455);
   U2326 : OAI22_X1 port map( A1 => n7739, A2 => n7740, B1 => n7986, B2 => 
                           n8615, ZN => n7989);
   U2330 : NAND2_X1 port map( A1 => n5433, A2 => n8423, ZN => n8422);
   U2349 : AOI21_X1 port map( B1 => n5432, B2 => n8349, A => n5434, ZN => n8424
                           );
   U2354 : OAI21_X1 port map( B1 => n6611, B2 => n6612, A => n6610, ZN => n6617
                           );
   U2356 : NAND3_X1 port map( A1 => n6837, A2 => n6833, A3 => n6834, ZN => 
                           n6994);
   U2390 : NAND2_X1 port map( A1 => n5543, A2 => n5542, ZN => n5568);
   U2448 : XNOR2_X1 port map( A => n6083, B => n6082, ZN => n7940);
   U2828 : XOR2_X1 port map( A => n5233, B => n5232, Z => n8430);
   U2936 : AOI21_X1 port map( B1 => n5498, B2 => n5497, A => n5496, ZN => n8431
                           );
   U3056 : AOI21_X1 port map( B1 => n5498, B2 => n5497, A => n5496, ZN => n5550
                           );
   U3086 : OR2_X1 port map( A1 => n5760, A2 => n5879, ZN => n8003);
   U3123 : XNOR2_X1 port map( A => n4999, B => n5102, ZN => n4351);
   U3266 : XNOR2_X1 port map( A => n4351, B => n4995, ZN => n5126);
   U3268 : BUF_X1 port map( A => n7080, Z => n4437);
   U3298 : NOR2_X1 port map( A1 => n7606, A2 => n8168, ZN => n8165);
   U3379 : BUF_X1 port map( A => n5845, Z => n8438);
   U3625 : NAND2_X1 port map( A1 => n5032, A2 => n5031, ZN => n8441);
   U3690 : OR2_X1 port map( A1 => n7489, A2 => n7488, ZN => n8443);
   U3796 : OR2_X2 port map( A1 => n4414, A2 => n8575, ZN => n8444);
   U3865 : BUF_X2 port map( A => n6388, Z => n8445);
   U4161 : AND2_X1 port map( A1 => n6629, A2 => n6628, ZN => n8448);
   U4162 : INV_X1 port map( A => n6089, ZN => n8449);
   U4176 : CLKBUF_X1 port map( A => n8115, Z => n8450);
   U4207 : OR2_X1 port map( A1 => n6719, A2 => n6720, ZN => n8451);
   U4245 : INV_X1 port map( A => n7065, ZN => n8452);
   U4309 : XOR2_X1 port map( A => n5115, B => n4405, Z => n8453);
   U4310 : INV_X1 port map( A => n4561, ZN => n8454);
   U4387 : INV_X1 port map( A => n4561, ZN => n6126);
   U4396 : INV_X1 port map( A => n6102, ZN => n8455);
   U4397 : AND2_X1 port map( A1 => n4808, A2 => n4809, ZN => n5794);
   U4437 : XOR2_X1 port map( A => n7019, B => n7115, Z => n8456);
   U4440 : OR2_X1 port map( A1 => n6713, A2 => n6712, ZN => n8458);
   U4533 : NAND2_X1 port map( A1 => n6738, A2 => n5879, ZN => n8004);
   U4586 : CLKBUF_X1 port map( A => n7929, Z => n8461);
   U4602 : AND2_X1 port map( A1 => n4550, A2 => n4549, ZN => n8462);
   U4623 : OR2_X1 port map( A1 => n6713, A2 => n6712, ZN => n6853);
   U4628 : BUF_X1 port map( A => n6988, Z => n8464);
   U4654 : OR2_X1 port map( A1 => n6909, A2 => n6908, ZN => n6988);
   U4661 : BUF_X1 port map( A => n6688, Z => n7323);
   U4690 : INV_X1 port map( A => n7594, ZN => n8466);
   U4691 : XOR2_X1 port map( A => n5551, B => n5553, Z => n5554);
   U4945 : NAND2_X1 port map( A1 => n6841, A2 => n6840, ZN => n8468);
   U5160 : NAND3_X1 port map( A1 => n5883, A2 => n5854, A3 => A_SIG_10_port, ZN
                           => n8469);
   U5164 : AND2_X1 port map( A1 => n6398, A2 => n6396, ZN => n8470);
   U5267 : OR2_X2 port map( A1 => n5937, A2 => n4514, ZN => n7254);
   U5274 : INV_X1 port map( A => n369, ZN => n8471);
   U5536 : BUF_X2 port map( A => n4963, Z => n7122);
   U5572 : AND2_X1 port map( A1 => n6783, A2 => n6782, ZN => n8472);
   U5631 : AND2_X1 port map( A1 => n8551, A2 => n6836, ZN => n8473);
   U5641 : NAND2_X1 port map( A1 => n6841, A2 => n6840, ZN => n8474);
   U5690 : AND2_X1 port map( A1 => n6922, A2 => n8451, ZN => n6970);
   U5693 : AOI21_X1 port map( B1 => n6054, B2 => n6055, A => n4365, ZN => n6077
                           );
   U5803 : XNOR2_X1 port map( A => n5820, B => n6055, ZN => n6074);
   U5805 : NOR2_X2 port map( A1 => n8186, A2 => n7600, ZN => n7625);
   U5809 : XOR2_X1 port map( A => n388, B => n8366, Z => n4658);
   U5810 : INV_X1 port map( A => n8530, ZN => n8479);
   U5811 : OR2_X1 port map( A1 => n8145, A2 => n8144, ZN => n8480);
   U5812 : OR2_X1 port map( A1 => n6465, A2 => n6464, ZN => n8481);
   U5816 : AND2_X1 port map( A1 => n7031, A2 => n7030, ZN => n8485);
   U5817 : AND2_X1 port map( A1 => n5882, A2 => n5881, ZN => n8487);
   U5818 : CLKBUF_X1 port map( A => n5168, Z => n4477);
   U5819 : BUF_X1 port map( A => n5396, Z => n8488);
   U5820 : NOR2_X1 port map( A1 => n4885, A2 => n8356, ZN => n5396);
   U5821 : XNOR2_X1 port map( A => n8489, B => n6525, ZN => n6223);
   U5823 : XOR2_X1 port map( A => n5826, B => n5825, Z => n8492);
   U5826 : XOR2_X1 port map( A => n8567, B => n5278, Z => n8495);
   U5827 : XOR2_X1 port map( A => n5548, B => n5547, Z => n8496);
   U5828 : CLKBUF_X1 port map( A => n5028, Z => n8497);
   U5829 : OR2_X1 port map( A1 => n6719, A2 => n6720, ZN => n6921);
   U5830 : OR2_X1 port map( A1 => n5869, A2 => n5868, ZN => n8498);
   U5832 : BUF_X1 port map( A => n7415, Z => n8500);
   U5833 : BUF_X1 port map( A => n7415, Z => n8501);
   U5834 : XOR2_X1 port map( A => n6359, B => n6592, Z => n8502);
   U5835 : INV_X1 port map( A => n8398, ZN => n8504);
   U5837 : INV_X1 port map( A => n8338, ZN => n8506);
   U5839 : INV_X1 port map( A => n5395, ZN => n8510);
   U5840 : INV_X1 port map( A => n4559, ZN => n6249);
   U5844 : CLKBUF_X1 port map( A => n6946, Z => n8513);
   U5845 : XNOR2_X1 port map( A => n382, B => n8360, ZN => n8514);
   U5846 : INV_X1 port map( A => n4560, ZN => n8515);
   U5847 : INV_X1 port map( A => n4560, ZN => n8516);
   U5848 : INV_X1 port map( A => n4560, ZN => n6248);
   U5849 : AOI21_X1 port map( B1 => n8025, B2 => n8026, A => n7923, ZN => n8517
                           );
   n8518 <= '0';
   n8520 <= '0';
   U5854 : NAND2_X1 port map( A1 => n8522, A2 => n8357, ZN => n6709);
   U5855 : NAND2_X1 port map( A1 => n6703, A2 => n359, ZN => n8522);
   U5856 : XNOR2_X1 port map( A => n5828, B => n5827, ZN => n4378);
   U5857 : NAND3_X1 port map( A1 => n4470, A2 => n4469, A3 => n4471, ZN => 
                           n5828);
   U2120 : NAND2_X2 port map( A1 => n6703, A2 => n8357, ZN => n4462);
   U2008 : AOI22_X2 port map( A1 => n6559, A2 => n6558, B1 => n6557, B2 => 
                           n6556, ZN => n4444);
   U1894 : OR2_X2 port map( A1 => n5760, A2 => n5879, ZN => n8434);
   U2117 : NAND3_X2 port map( A1 => n4432, A2 => n7733, A3 => n8443, ZN => 
                           n4459);
   U5264 : AOI21_X2 port map( B1 => n8121, B2 => n7725, A => n7724, ZN => n7983
                           );
   U1890 : BUF_X2 port map( A => n6342, Z => n7439);
   U2161 : BUF_X2 port map( A => n6889, Z => n4490);
   U1790 : NOR2_X2 port map( A1 => n6367, A2 => n6366, ZN => n6395);
   U2462 : OAI22_X2 port map( A1 => n6381, A2 => n6252, B1 => n6382, B2 => 
                           n6251, ZN => n8429);
   U1832 : OR2_X2 port map( A1 => n6544, A2 => n6547, ZN => n6490);
   U1801 : BUF_X2 port map( A => n4817, Z => n6251);
   U1776 : NAND2_X2 port map( A1 => n6343, A2 => n5272, ZN => n6800);
   U2223 : OR2_X1 port map( A1 => n7152, A2 => n7151, ZN => n7278);
   U2970 : NOR2_X1 port map( A1 => n8353, A2 => n384, ZN => n6227);
   U2052 : OR2_X1 port map( A1 => n5910, A2 => n5909, ZN => n6211);
   I1_B_SIG_reg_3_inst : DFF_X1 port map( D => FP_B(3), CK => clk, Q => n8328, 
                           QN => n386);
   I3_SIG_out_round_reg_26_U4 : MUX2_X1 port map( A => n8375, B => n4527, S => 
                           n8404, Z => n8608);
   I3_SIG_out_round_reg_26_inst : DFF_X1 port map( D => n8608, CK => clk, Q => 
                           SIG_out_round_26_port, QN => n_1149);
   I2_prod_tmp_reg_38_inst : DFFRS_X1 port map( D => I2_dtemp_38_port, CK => 
                           clk, RN => n8607, SN => n8607, Q => 
                           I2_SIG_in_int_18_port, QN => n_1150);
   I1_B_SIG_reg_20_inst : DFF_X2 port map( D => FP_B(20), CK => clk, Q => n8349
                           , QN => n8423);
   I2_prod_tmp_reg_44_inst : DFFRS_X1 port map( D => I2_dtemp_44_port, CK => 
                           clk, RN => n8606, SN => n8606, Q => 
                           I2_SIG_in_int_24_port, QN => n_1151);
   I1_B_SIG_reg_18_inst : DFF_X1 port map( D => FP_B(18), CK => clk, Q => n8329
                           , QN => n363);
   I1_B_SIG_reg_6_inst : DFF_X1 port map( D => FP_B(6), CK => clk, Q => n8352, 
                           QN => n390);
   I2_prod_tmp_reg_40_inst : DFF_X1 port map( D => I2_dtemp_40_port, CK => clk,
                           Q => I2_SIG_in_int_20_port, QN => n_1152);
   I2_prod_tmp_reg_39_inst : DFF_X1 port map( D => I2_dtemp_39_port, CK => clk,
                           Q => I2_SIG_in_int_19_port, QN => n_1153);
   U2401 : BUF_X1 port map( A => n385, Z => n4892);
   U2360 : BUF_X1 port map( A => n394, Z => n4961);
   I1_B_SIG_reg_12_inst : DFF_X1 port map( D => FP_B(12), CK => clk, Q => n4381
                           , QN => n373);
   U2350 : BUF_X2 port map( A => n382, Z => n5883);
   U1736 : BUF_X1 port map( A => n8338, Z => n5854);
   U1805 : NAND2_X1 port map( A1 => n8358, A2 => n8395, ZN => n7947);
   U1905 : BUF_X1 port map( A => A_SIG_16_port, Z => n6706);
   U1803 : CLKBUF_X2 port map( A => n388, Z => n6244);
   U1889 : BUF_X1 port map( A => n5866, Z => n8476);
   U1729 : BUF_X1 port map( A => n6688, Z => n8465);
   U2341 : BUF_X1 port map( A => n376, Z => n6606);
   U2066 : BUF_X1 port map( A => n7195, Z => n4487);
   U1880 : BUF_X1 port map( A => n7254, Z => n7773);
   U1856 : AND2_X1 port map( A1 => n5989, A2 => n5988, ZN => n6171);
   I2_prod_tmp_reg_28_inst : DFF_X1 port map( D => I2_dtemp_28_port, CK => clk,
                           Q => I2_SIG_in_int_8_port, QN => n_1154);
   I2_prod_tmp_reg_30_inst : DFF_X1 port map( D => I2_dtemp_30_port, CK => clk,
                           Q => I2_SIG_in_int_10_port, QN => n_1155);
   I2_prod_tmp_reg_26_inst : DFF_X1 port map( D => I2_dtemp_26_port, CK => clk,
                           Q => I2_SIG_in_int_6_port, QN => n_1156);
   I2_prod_tmp_reg_32_inst : DFF_X1 port map( D => n8405, CK => clk, Q => 
                           I2_SIG_in_int_12_port, QN => n_1157);
   I2_prod_tmp_reg_47_inst : DFF_X1 port map( D => n8367, CK => clk, Q => 
                           I2_SIG_in_int_27_port, QN => n_1158);
   I1_B_SIG_reg_7_inst : DFF_X2 port map( D => FP_B(7), CK => clk, Q => n8333, 
                           QN => n362);
   I1_B_SIG_reg_15_inst : DFF_X2 port map( D => FP_B(15), CK => clk, Q => n8332
                           , QN => n377);
   U1739 : OR2_X1 port map( A1 => n7583, A2 => n8624, ZN => n7593);
   U1743 : AND2_X1 port map( A1 => n7987, A2 => n8613, ZN => n8612);
   U1745 : AND2_X1 port map( A1 => n5907, A2 => n5951, ZN => n6199);
   U1748 : NAND2_X1 port map( A1 => n8621, A2 => n8620, ZN => n5894);
   U1750 : BUF_X2 port map( A => SIG_in_27_port, Z => n8089);
   U1751 : NAND2_X1 port map( A1 => n5921, A2 => n8487, ZN => n8620);
   U1755 : BUF_X1 port map( A => n8478, Z => n8596);
   U1757 : OR2_X1 port map( A1 => n6692, A2 => n6691, ZN => n6839);
   U1758 : BUF_X2 port map( A => n5051, Z => n7861);
   U1760 : BUF_X2 port map( A => n6343, Z => n6593);
   U1763 : BUF_X1 port map( A => n4559, Z => n5395);
   U1765 : BUF_X1 port map( A => n4632, Z => n7051);
   U1766 : CLKBUF_X2 port map( A => n393, Z => n6343);
   U1767 : BUF_X1 port map( A => n6705, Z => n6363);
   U1768 : CLKBUF_X1 port map( A => n4885, Z => n5055);
   U1788 : CLKBUF_X1 port map( A => n5844, Z => n8436);
   U1791 : CLKBUF_X1 port map( A => n4808, Z => n5846);
   U1792 : AOI21_X1 port map( B1 => n6306, B2 => n6307, A => n6305, ZN => n6310
                           );
   U1793 : NAND2_X1 port map( A1 => n5385, A2 => n5777, ZN => n8559);
   U1802 : BUF_X1 port map( A => n7080, Z => n7325);
   U1804 : OR2_X1 port map( A1 => n6351, A2 => n6350, ZN => n6620);
   U1806 : NAND2_X1 port map( A1 => n6127, A2 => n8510, ZN => n6284);
   U1810 : CLKBUF_X1 port map( A => n5040, Z => n5041);
   U1811 : AOI22_X1 port map( A1 => n6429, A2 => n4375, B1 => n6428, B2 => 
                           n6427, ZN => n6436);
   U1812 : OAI21_X1 port map( B1 => n6586, B2 => n6585, A => n6584, ZN => n8587
                           );
   U1814 : NAND2_X1 port map( A1 => n5385, A2 => n5777, ZN => n7090);
   U1815 : BUF_X1 port map( A => n7086, Z => n7665);
   U1822 : BUF_X1 port map( A => B_SIG_8_port, Z => n7945);
   U1824 : BUF_X1 port map( A => n4963, Z => n6812);
   U1829 : INV_X1 port map( A => n6331, ZN => n8625);
   U1830 : OR2_X1 port map( A1 => n6238, A2 => n6239, ZN => n6437);
   U1831 : BUF_X1 port map( A => n364, Z => n7506);
   U1849 : AND2_X1 port map( A1 => n7129, A2 => n7130, ZN => n7174);
   U1853 : OR2_X1 port map( A1 => n7302, A2 => n7301, ZN => n7401);
   U1862 : XNOR2_X1 port map( A => n8626, B => n8625, ZN => n6338);
   U1863 : CLKBUF_X1 port map( A => n6974, Z => n6945);
   U1865 : XNOR2_X1 port map( A => n6242, B => n6440, ZN => n6445);
   U1866 : BUF_X1 port map( A => n364, Z => n7769);
   U1869 : CLKBUF_X1 port map( A => n7599, Z => n7613);
   U1870 : CLKBUF_X1 port map( A => n7635, Z => n4483);
   U1876 : CLKBUF_X1 port map( A => n6517, Z => n6214);
   U1882 : CLKBUF_X1 port map( A => n5861, Z => n7087);
   U1884 : CLKBUF_X1 port map( A => n7161, Z => n7167);
   U1893 : CLKBUF_X1 port map( A => n6546, Z => n6512);
   U1900 : OR2_X1 port map( A1 => n6517, A2 => n6516, ZN => n6541);
   U1902 : NOR2_X1 port map( A1 => n8615, A2 => n8614, ZN => n8613);
   U1903 : AND3_X1 port map( A1 => n8208, A2 => n7587, A3 => n8207, ZN => n7585
                           );
   U1908 : CLKBUF_X1 port map( A => n7629, Z => n7959);
   U1913 : CLKBUF_X1 port map( A => n8033, Z => n4463);
   U1927 : CLKBUF_X1 port map( A => n7727, Z => n4399);
   U1928 : CLKBUF_X1 port map( A => n8089, Z => n8279);
   U1931 : NAND2_X1 port map( A1 => n8126, A2 => n8129, ZN => n8526);
   U1933 : OR2_X1 port map( A1 => n7650, A2 => n7483, ZN => n8527);
   U1936 : OR2_X1 port map( A1 => n7650, A2 => n7483, ZN => n7733);
   U1948 : INV_X1 port map( A => n7253, ZN => n8528);
   U1955 : NAND2_X1 port map( A1 => n7364, A2 => n7365, ZN => n8529);
   U1960 : BUF_X1 port map( A => n4632, Z => n7084);
   U1967 : INV_X1 port map( A => n6811, ZN => n8530);
   U1971 : BUF_X1 port map( A => n5030, Z => n6811);
   U1975 : CLKBUF_X1 port map( A => n7940, Z => n8428);
   U1986 : NAND2_X1 port map( A1 => n4461, A2 => n8362, ZN => n8610);
   U2005 : NAND2_X1 port map( A1 => n6031, A2 => n6029, ZN => n8531);
   U2010 : NAND2_X1 port map( A1 => n6060, A2 => n6059, ZN => n8532);
   U2011 : NAND2_X1 port map( A1 => n5276, A2 => n5275, ZN => n8533);
   U2012 : CLKBUF_X1 port map( A => n6558, Z => n8534);
   U2019 : INV_X1 port map( A => n5395, ZN => n8535);
   U2025 : OR2_X1 port map( A1 => n7963, A2 => n8618, ZN => n7964);
   U2034 : AND2_X2 port map( A1 => n4364, A2 => n6259, ZN => n4560);
   U2036 : AND2_X2 port map( A1 => n6787, A2 => n6786, ZN => n7022);
   U2037 : OR2_X1 port map( A1 => n6665, A2 => n6664, ZN => n8628);
   U2044 : CLKBUF_X1 port map( A => n7493, Z => n8578);
   U2046 : NAND2_X2 port map( A1 => n6738, A2 => n5879, ZN => n8459);
   U2050 : NAND2_X2 port map( A1 => n5837, A2 => n5836, ZN => n6153);
   U2057 : CLKBUF_X1 port map( A => n6681, Z => n8536);
   U2077 : CLKBUF_X1 port map( A => n5149, Z => n8537);
   U2081 : CLKBUF_X1 port map( A => n8355, Z => n8538);
   U2121 : OAI211_X1 port map( C1 => n5685, C2 => n5490, A => n5670, B => n5489
                           , ZN => n8539);
   U2124 : OR2_X1 port map( A1 => n5147, A2 => n5146, ZN => n5205);
   U2127 : XNOR2_X1 port map( A => n5820, B => n6055, ZN => n8540);
   U2134 : AND2_X1 port map( A1 => n8529, A2 => n8129, ZN => n8541);
   U2138 : INV_X1 port map( A => n7488, ZN => n8542);
   U2142 : NAND2_X1 port map( A1 => n8086, A2 => n6561, ZN => n8484);
   U2143 : CLKBUF_X1 port map( A => n5744, Z => n5749);
   U2152 : INV_X1 port map( A => n7690, ZN => n7771);
   U2155 : XNOR2_X1 port map( A => n6152, B => n6153, ZN => n8543);
   U2156 : XNOR2_X1 port map( A => n5645, B => n5968, ZN => n8544);
   U2175 : CLKBUF_X1 port map( A => n8129, Z => n4426);
   U2212 : OAI211_X1 port map( C1 => n6582, C2 => n6581, A => n6580, B => n6579
                           , ZN => n8545);
   U2215 : CLKBUF_X1 port map( A => n5844, Z => n8546);
   U2226 : CLKBUF_X1 port map( A => n8103, Z => n8104);
   U2235 : CLKBUF_X1 port map( A => n5845, Z => n8547);
   U2255 : INV_X1 port map( A => n7253, ZN => n7499);
   U2263 : CLKBUF_X1 port map( A => n7602, Z => n8147);
   U2300 : XOR2_X1 port map( A => n6265, B => n6434, Z => n8548);
   U2301 : AOI22_X2 port map( A1 => n5644, A2 => n5643, B1 => n5642, B2 => 
                           n5641, ZN => n5968);
   U2319 : CLKBUF_X1 port map( A => n7723, Z => n8229);
   U2334 : AND2_X1 port map( A1 => n6250, A2 => n6251, ZN => n8549);
   U2362 : XNOR2_X1 port map( A => n7019, B => n8603, ZN => n8550);
   U2446 : XOR2_X1 port map( A => n6806, B => n7027, Z => n8551);
   U2567 : AOI22_X2 port map( A1 => n7282, A2 => n7281, B1 => n7280, B2 => 
                           n7289, ZN => n7607);
   U2598 : BUF_X1 port map( A => n5793, Z => n8552);
   U2711 : BUF_X1 port map( A => n5793, Z => n8553);
   U2818 : NOR2_X1 port map( A1 => n4810, A2 => n4809, ZN => n5793);
   U2823 : CLKBUF_X1 port map( A => n384, Z => n5620);
   U2846 : XNOR2_X1 port map( A => n6816, B => n6882, ZN => n8554);
   U2862 : XNOR2_X1 port map( A => n6928, B => n6927, ZN => n8555);
   U2946 : OAI211_X1 port map( C1 => n7227, C2 => n386, A => n5647, B => n4530,
                           ZN => n8556);
   U2969 : BUF_X1 port map( A => n6028, Z => n8557);
   U2979 : NAND2_X1 port map( A1 => n8077, A2 => n4444, ZN => n8558);
   U3065 : AND2_X2 port map( A1 => n8040, A2 => n8042, ZN => n7943);
   U3087 : AOI22_X2 port map( A1 => n5451, A2 => n5450, B1 => n5449, B2 => 
                           n5448, ZN => n5586);
   U3127 : NAND2_X2 port map( A1 => n6032, A2 => n6031, ZN => n6521);
   U3288 : NAND2_X1 port map( A1 => n6597, A2 => n6596, ZN => n8560);
   U3375 : NAND2_X1 port map( A1 => n4459, A2 => n7495, ZN => n8561);
   U3376 : XOR2_X1 port map( A => n7575, B => n7574, Z => n8562);
   U3382 : OAI22_X1 port map( A1 => n7986, A2 => n8615, B1 => n7740, B2 => 
                           n7739, ZN => n8563);
   U3430 : CLKBUF_X1 port map( A => n8057, Z => n8075);
   U3452 : CLKBUF_X1 port map( A => n390, Z => n8564);
   U3578 : AOI22_X1 port map( A1 => n6434, A2 => n6433, B1 => n8415, B2 => 
                           n6431, ZN => n8565);
   U3582 : CLKBUF_X1 port map( A => n6493, Z => n8566);
   U3636 : XNOR2_X1 port map( A => n6441, B => n6653, ZN => n6493);
   U3637 : OAI211_X1 port map( C1 => n6404, C2 => n6403, A => n6402, B => n6401
                           , ZN => n6647);
   U3673 : AND2_X1 port map( A1 => n8339, A2 => n365, ZN => n5302);
   U3692 : CLKBUF_X1 port map( A => n5572, Z => n5570);
   U3701 : CLKBUF_X1 port map( A => n6528, Z => n6502);
   U3717 : XNOR2_X1 port map( A => n8533, B => n5481, ZN => n8567);
   U3747 : AND2_X1 port map( A1 => n4445, A2 => n7796, ZN => n8627);
   U3786 : CLKBUF_X1 port map( A => n7227, Z => n8568);
   U3830 : NAND2_X1 port map( A1 => n6093, A2 => n6091, ZN => n8569);
   U3841 : XNOR2_X1 port map( A => n5494, B => n5669, ZN => n8570);
   U3858 : XNOR2_X1 port map( A => n6496, B => n6495, ZN => n8571);
   U3863 : XOR2_X1 port map( A => n8543, B => n6149, Z => n8572);
   U3907 : AND2_X1 port map( A1 => n6139, A2 => n6138, ZN => n8573);
   U3914 : XOR2_X1 port map( A => n8571, B => n6497, Z => n8574);
   U3983 : NOR2_X1 port map( A1 => n6223, A2 => n6224, ZN => n8575);
   U3999 : CLKBUF_X1 port map( A => n6342, Z => n7508);
   U4000 : XNOR2_X1 port map( A => n6752, B => n6858, ZN => n8576);
   U4001 : XNOR2_X1 port map( A => n6752, B => n6858, ZN => n6933);
   U4003 : BUF_X2 port map( A => n4632, Z => n8577);
   U4012 : CLKBUF_X1 port map( A => n6911, Z => n8579);
   U4047 : NAND2_X1 port map( A1 => n6703, A2 => n8357, ZN => n4461);
   U4055 : CLKBUF_X1 port map( A => n8157, Z => n8580);
   U4117 : CLKBUF_X1 port map( A => n6696, Z => n8581);
   U4139 : BUF_X2 port map( A => n6696, Z => n8582);
   U4184 : XNOR2_X1 port map( A => n5401, B => n5597, ZN => n8583);
   U4226 : CLKBUF_X1 port map( A => n7492, Z => n8584);
   U4234 : NOR2_X1 port map( A1 => n7605, A2 => n4441, ZN => n8585);
   U4238 : NOR2_X1 port map( A1 => n7605, A2 => n4441, ZN => n7479);
   U4251 : CLKBUF_X1 port map( A => n8558, Z => n8586);
   U4257 : OAI21_X1 port map( B1 => n6586, B2 => n6585, A => n6584, ZN => n4416
                           );
   U4274 : XNOR2_X2 port map( A => n6554, B => n6553, ZN => n8077);
   U4423 : CLKBUF_X1 port map( A => n7605, Z => n7606);
   U4472 : CLKBUF_X1 port map( A => n6863, Z => n8588);
   U4474 : XNOR2_X1 port map( A => n6862, B => n6863, ZN => n8589);
   U4500 : AND2_X1 port map( A1 => n8057, A2 => n8586, ZN => n8590);
   U4530 : AOI22_X1 port map( A1 => n6172, A2 => n6171, B1 => n6170, B2 => 
                           n6169, ZN => n8591);
   U4597 : XNOR2_X1 port map( A => n7267, B => n7349, ZN => n8592);
   U4621 : NAND2_X1 port map( A1 => n4961, A2 => n8629, ZN => n8593);
   U4637 : NAND2_X1 port map( A1 => n4961, A2 => n8629, ZN => n7123);
   U4745 : AND2_X1 port map( A1 => n8471, A2 => n8340, ZN => n8629);
   U4746 : AND2_X2 port map( A1 => n5161, A2 => n5160, ZN => n5168);
   U4747 : CLKBUF_X1 port map( A => n7378, Z => n7608);
   U4758 : OAI21_X2 port map( B1 => n5441, B2 => n5501, A => n5500, ZN => n5584
                           );
   U4840 : OR2_X2 port map( A1 => n6911, A2 => n6910, ZN => n6935);
   U4854 : MUX2_X1 port map( A => n8593, B => n6812, S => n360, Z => n6608);
   U4877 : AND2_X2 port map( A1 => n4993, A2 => n8369, ZN => n5226);
   U4938 : INV_X1 port map( A => n6562, ZN => n8594);
   U5049 : XNOR2_X1 port map( A => n6488, B => n6670, ZN => n8086);
   U5055 : OR2_X1 port map( A1 => n7650, A2 => n7651, ZN => n8096);
   U5059 : AOI21_X2 port map( B1 => n7629, B2 => n7643, A => n7498, ZN => n8208
                           );
   U5061 : NOR2_X2 port map( A1 => n7729, A2 => n8212, ZN => n7986);
   U5064 : BUF_X1 port map( A => n8478, Z => n8595);
   U5101 : NAND2_X1 port map( A1 => n4544, A2 => n8366, ZN => n8478);
   U5140 : AOI21_X1 port map( B1 => n8025, B2 => n8026, A => n7923, ZN => n8597
                           );
   U5141 : AOI22_X1 port map( A1 => n4456, A2 => n6936, B1 => n6935, B2 => 
                           n6934, ZN => n8598);
   U5142 : OAI22_X1 port map( A1 => n4518, A2 => n6587, B1 => n6592, B2 => 
                           n6589, ZN => n8599);
   U5195 : CLKBUF_X1 port map( A => n4421, Z => n8600);
   U5270 : NOR2_X1 port map( A1 => n7721, A2 => n8096, ZN => n8601);
   U5529 : NOR2_X1 port map( A1 => n7721, A2 => n8096, ZN => n4412);
   U5535 : XNOR2_X1 port map( A => n7063, B => n7153, ZN => n8602);
   U5548 : XNOR2_X1 port map( A => n7018, B => n7144, ZN => n8603);
   U5550 : XOR2_X1 port map( A => n8550, B => n7075, Z => n8604);
   U5552 : NAND2_X1 port map( A1 => n4459, A2 => n7495, ZN => n8605);
   n8606 <= '1';
   n8607 <= '1';
   U5806 : NAND2_X1 port map( A1 => n8610, A2 => n8609, ZN => n5840);
   U5807 : NAND2_X1 port map( A1 => n7054, A2 => n7945, ZN => n8609);
   U5808 : NAND2_X4 port map( A1 => n4993, A2 => n8369, ZN => n7324);
   U5813 : AND2_X2 port map( A1 => n358, A2 => n394, ZN => n4993);
   U5814 : OR2_X1 port map( A1 => n6380, A2 => n6379, ZN => n6407);
   U5815 : OAI211_X1 port map( C1 => n7994, C2 => n7995, A => n8611, B => n7992
                           , ZN => n8411);
   U5822 : NAND2_X1 port map( A1 => n7995, A2 => n8612, ZN => n8611);
   U5824 : INV_X1 port map( A => n7994, ZN => n8614);
   U5825 : INV_X1 port map( A => n7988, ZN => n8615);
   U5831 : OR2_X1 port map( A1 => n7140, A2 => n7141, ZN => n7188);
   U5836 : OR2_X1 port map( A1 => n4461, A2 => n8392, ZN => n8632);
   U5838 : OAI21_X1 port map( B1 => n6292, B2 => n6293, A => n6291, ZN => n6295
                           );
   U5841 : OR2_X1 port map( A1 => n8555, A2 => n7365, ZN => n7601);
   U5842 : AND2_X2 port map( A1 => n6287, A2 => n6286, ZN => n6292);
   U5843 : XNOR2_X1 port map( A => n8617, B => n8616, ZN => n8489);
   U5851 : INV_X1 port map( A => n6524, ZN => n8616);
   U5853 : NAND2_X1 port map( A1 => n6096, A2 => n6095, ZN => n8617);
   U5858 : NAND2_X1 port map( A1 => n7960, A2 => n8619, ZN => n8618);
   U5859 : INV_X1 port map( A => n7962, ZN => n8619);
   U5860 : INV_X1 port map( A => n5894, ZN => n5893);
   U5861 : NAND2_X1 port map( A1 => n5889, A2 => n5918, ZN => n8621);
   U5862 : NOR2_X1 port map( A1 => n8622, A2 => n7011, ZN => n7015);
   U5863 : NAND2_X1 port map( A1 => n7013, A2 => n8623, ZN => n8622);
   U5864 : NAND2_X1 port map( A1 => n7012, A2 => n8331, ZN => n8623);
   U5865 : INV_X1 port map( A => n7585, ZN => n8624);
   U5866 : NAND2_X1 port map( A1 => n6330, A2 => n6329, ZN => n8626);
   U5867 : NAND2_X1 port map( A1 => n4450, A2 => n7368, ZN => n8103);
   U5868 : XNOR2_X1 port map( A => n4475, B => n4474, ZN => n7368);
   U5869 : NAND2_X1 port map( A1 => n4449, A2 => n8627, ZN => n4347);
   U5870 : NAND3_X1 port map( A1 => n6663, A2 => n6662, A3 => n8628, ZN => 
                           n4429);
   U5871 : AND2_X2 port map( A1 => n8353, A2 => n5620, ZN => n6703);
   U5872 : XNOR2_X1 port map( A => n8630, B => n6939, ZN => n6967);
   U5873 : XNOR2_X1 port map( A => n6971, B => n6938, ZN => n8630);
   U5874 : NAND2_X1 port map( A1 => n8632, A2 => n8631, ZN => n6367);
   U5875 : NAND2_X1 port map( A1 => n6361, A2 => n8392, ZN => n8631);

end SYN_pipeline;
