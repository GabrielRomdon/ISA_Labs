
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_FPmul is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_FPmul;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_20 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_20;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_19 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_19;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_18 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_18;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_17 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_17;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_16 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_16;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_15 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_15;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_13 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_13;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_22 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_22;

architecture SYN_STRUCTURAL of RCA_generic_N2_22 is

   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102698, n_1002 : std_logic;

begin
   
   net102698 <= '0';
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => net102698, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1002);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_20 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_20;

architecture SYN_STRUCTURAL of RCA_generic_N2_20 is

   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102698, n_1005 : std_logic;

begin
   
   net102698 <= '0';
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => net102698, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1005);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_21 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_21;

architecture SYN_STRUCTURAL of RCA_generic_N2_21 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102701, n_1008 : std_logic;

begin
   
   net102701 <= '0';
   FAI_1 : FA_42 port map( A => A(0), B => B(0), Ci => net102701, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_41 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1008);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_19 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_19;

architecture SYN_STRUCTURAL of RCA_generic_N2_19 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102701, n_1011 : std_logic;

begin
   
   net102701 <= '0';
   FAI_1 : FA_38 port map( A => A(0), B => B(0), Ci => net102701, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_37 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1011);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_68 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_68;

architecture SYN_BEHAVIORAL of PG_GENERAL_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_76 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_76;

architecture SYN_BEHAVIORAL of PG_GENERAL_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_75 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_75;

architecture SYN_BEHAVIORAL of PG_GENERAL_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_71 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_71;

architecture SYN_BEHAVIORAL of PG_GENERAL_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_69 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_69;

architecture SYN_BEHAVIORAL of PG_GENERAL_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_79 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_79;

architecture SYN_BEHAVIORAL of PG_GENERAL_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_78 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_78;

architecture SYN_BEHAVIORAL of PG_GENERAL_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_73 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_73;

architecture SYN_BEHAVIORAL of PG_GENERAL_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_49 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_49;

architecture SYN_BEHAVIORAL of PG_GENERAL_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_48 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_48;

architecture SYN_BEHAVIORAL of PG_GENERAL_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_47 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_47;

architecture SYN_BEHAVIORAL of PG_GENERAL_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_46 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_46;

architecture SYN_BEHAVIORAL of PG_GENERAL_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_45 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_45;

architecture SYN_BEHAVIORAL of PG_GENERAL_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_40 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_40;

architecture SYN_BEHAVIORAL of PG_GENERAL_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_33 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_33;

architecture SYN_BEHAVIORAL of PG_GENERAL_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_30 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_30;

architecture SYN_BEHAVIORAL of PG_GENERAL_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_28 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_28;

architecture SYN_BEHAVIORAL of PG_GENERAL_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_26 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_26;

architecture SYN_BEHAVIORAL of PG_GENERAL_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_18 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_18;

architecture SYN_BEHAVIORAL of PG_GENERAL_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_13 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_13;

architecture SYN_BEHAVIORAL of G_GENERAL_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_48 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_48;

architecture SYN_BEHAVIORAL of PG_NET_48 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_47 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_47;

architecture SYN_BEHAVIORAL of PG_NET_47 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_43 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_43;

architecture SYN_BEHAVIORAL of PG_NET_43 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_41 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_41;

architecture SYN_BEHAVIORAL of PG_NET_41 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_40 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_40;

architecture SYN_BEHAVIORAL of PG_NET_40 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_46 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_46;

architecture SYN_BEHAVIORAL of PG_NET_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_34 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_34;

architecture SYN_BEHAVIORAL of PG_NET_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_36 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_36;

architecture SYN_BEHAVIORAL of PG_NET_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_30 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_30;

architecture SYN_BEHAVIORAL of PG_NET_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_28 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_28;

architecture SYN_BEHAVIORAL of PG_NET_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_22 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_22;

architecture SYN_BEHAVIORAL of PG_NET_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_33 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_33;

architecture SYN_BEHAVIORAL of PG_NET_33 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : INV_X1 port map( A => B, ZN => n1);
   U3 : XNOR2_X1 port map( A => A, B => n1, ZN => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_21 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_21;

architecture SYN_BEHAVIORAL of PG_NET_21 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : INV_X1 port map( A => B, ZN => n1);
   U3 : XNOR2_X1 port map( A => A, B => n1, ZN => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_24 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_24;

architecture SYN_BEHAVIORAL of PG_NET_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_23 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_23;

architecture SYN_BEHAVIORAL of PG_NET_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_61 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_61;

architecture SYN_BEHAVIORAL of PG_NET_61 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_57 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_57;

architecture SYN_BEHAVIORAL of PG_NET_57 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_56 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_56;

architecture SYN_BEHAVIORAL of PG_NET_56 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_55 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_55;

architecture SYN_BEHAVIORAL of PG_NET_55 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_51 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_51;

architecture SYN_BEHAVIORAL of PG_NET_51 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_39 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_39;

architecture SYN_BEHAVIORAL of PG_NET_39 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_20 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_20;

architecture SYN_BEHAVIORAL of PG_NET_20 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_568 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_568;

architecture SYN_BEHAVIORAL of FA_568 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_561 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_561;

architecture SYN_BEHAVIORAL of FA_561 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U5 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_586 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_586;

architecture SYN_BEHAVIORAL of FA_586 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_548 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_548;

architecture SYN_BEHAVIORAL of FA_548 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_564 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_564;

architecture SYN_BEHAVIORAL of FA_564 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_481;

architecture SYN_BEHAVIORAL of FA_481 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_463;

architecture SYN_BEHAVIORAL of FA_463 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_575 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_575;

architecture SYN_BEHAVIORAL of FA_575 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_507;

architecture SYN_BEHAVIORAL of FA_507 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_461;

architecture SYN_BEHAVIORAL of FA_461 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_517 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_517;

architecture SYN_BEHAVIORAL of FA_517 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_464;

architecture SYN_BEHAVIORAL of FA_464 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_531 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_531;

architecture SYN_BEHAVIORAL of FA_531 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_530 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_530;

architecture SYN_BEHAVIORAL of FA_530 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_516 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_516;

architecture SYN_BEHAVIORAL of FA_516 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_415;

architecture SYN_BEHAVIORAL of FA_415 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_377;

architecture SYN_BEHAVIORAL of FA_377 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_337;

architecture SYN_BEHAVIORAL of FA_337 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_502;

architecture SYN_BEHAVIORAL of FA_502 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_504;

architecture SYN_BEHAVIORAL of FA_504 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_545 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_545;

architecture SYN_BEHAVIORAL of FA_545 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_533 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_533;

architecture SYN_BEHAVIORAL of FA_533 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_532 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_532;

architecture SYN_BEHAVIORAL of FA_532 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_503;

architecture SYN_BEHAVIORAL of FA_503 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_484;

architecture SYN_BEHAVIORAL of FA_484 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_480 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_480;

architecture SYN_BEHAVIORAL of FA_480 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_477 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_477;

architecture SYN_BEHAVIORAL of FA_477 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_459;

architecture SYN_BEHAVIORAL of FA_459 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_410;

architecture SYN_BEHAVIORAL of FA_410 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_354 is

   port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_354;

architecture SYN_BEHAVIORAL of FA_354 is

begin
   S_BAR <= A_BAR;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_353 is

   port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_353;

architecture SYN_BEHAVIORAL of FA_353 is

begin
   S_BAR <= A_BAR;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_352 is

   port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_352;

architecture SYN_BEHAVIORAL of FA_352 is

begin
   S_BAR <= A_BAR;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL_architecture of FA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL_architecture of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_29 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_29;

architecture SYN_STRUCTURAL of RCA_generic_N2_29 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102703, n_1055 : std_logic;

begin
   
   net102703 <= '0';
   FAI_1 : FA_58 port map( A => A(0), B => B(0), Ci => net102703, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_57 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1055);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_542 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_542;

architecture SYN_BEHAVIORAL of FA_542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_540 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_540;

architecture SYN_BEHAVIORAL of FA_540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_489 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_489;

architecture SYN_BEHAVIORAL of FA_489 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_488 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_488;

architecture SYN_BEHAVIORAL of FA_488 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_487 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_487;

architecture SYN_BEHAVIORAL of FA_487 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_413;

architecture SYN_BEHAVIORAL of FA_413 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_515 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_515;

architecture SYN_BEHAVIORAL of FA_515 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_514 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_514;

architecture SYN_BEHAVIORAL of FA_514 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_513 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_513;

architecture SYN_BEHAVIORAL of FA_513 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_512 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_512;

architecture SYN_BEHAVIORAL of FA_512 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_505;

architecture SYN_BEHAVIORAL of FA_505 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_485 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_485;

architecture SYN_BEHAVIORAL of FA_485 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_417;

architecture SYN_BEHAVIORAL of FA_417 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_416;

architecture SYN_BEHAVIORAL of FA_416 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_380;

architecture SYN_BEHAVIORAL of FA_380 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_379;

architecture SYN_BEHAVIORAL of FA_379 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_378 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_378;

architecture SYN_BEHAVIORAL of FA_378 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_376;

architecture SYN_BEHAVIORAL of FA_376 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_375;

architecture SYN_BEHAVIORAL of FA_375 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_344;

architecture SYN_BEHAVIORAL of FA_344 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  Co, S : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  Co, S : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  Co, S : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_420;

architecture SYN_BEHAVIORAL of FA_420 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_419;

architecture SYN_BEHAVIORAL of FA_419 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_418;

architecture SYN_BEHAVIORAL of FA_418 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_373;

architecture SYN_BEHAVIORAL of FA_373 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_343;

architecture SYN_BEHAVIORAL of FA_343 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL_architecture of FA_42 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL_architecture of FA_38 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_41 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_41;

architecture SYN_rtl of HA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_40 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_40;

architecture SYN_rtl of HA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_39 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_39;

architecture SYN_rtl of HA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_38 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_38;

architecture SYN_rtl of HA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_37 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_37;

architecture SYN_rtl of HA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_36 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_36;

architecture SYN_rtl of HA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_35 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_35;

architecture SYN_rtl of HA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_34 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_34;

architecture SYN_rtl of HA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_32 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_32;

architecture SYN_rtl of HA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_31 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_31;

architecture SYN_rtl of HA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_29 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_29;

architecture SYN_rtl of HA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_28 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_28;

architecture SYN_rtl of HA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_26 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_26;

architecture SYN_rtl of HA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_25 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_25;

architecture SYN_rtl of HA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_24 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_24;

architecture SYN_rtl of HA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_23 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_23;

architecture SYN_rtl of HA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_20 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_20;

architecture SYN_rtl of HA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_19 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_19;

architecture SYN_rtl of HA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_17 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_17;

architecture SYN_rtl of HA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_16 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_16;

architecture SYN_rtl of HA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_14 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_14;

architecture SYN_rtl of HA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_13 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_13;

architecture SYN_rtl of HA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_10 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_10;

architecture SYN_rtl of HA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_8 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_8;

architecture SYN_rtl of HA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_7 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_7;

architecture SYN_rtl of HA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_5 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_5;

architecture SYN_rtl of HA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_4 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_4;

architecture SYN_rtl of HA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_2 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_2;

architecture SYN_rtl of HA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_1 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_1;

architecture SYN_rtl of HA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_22 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_22;

architecture SYN_BEHAVIORAL of G_GENERAL_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_20 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_20;

architecture SYN_BEHAVIORAL of G_GENERAL_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_19 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_19;

architecture SYN_BEHAVIORAL of G_GENERAL_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_18 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_18;

architecture SYN_BEHAVIORAL of G_GENERAL_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_16 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_16;

architecture SYN_BEHAVIORAL of G_GENERAL_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_15 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_15;

architecture SYN_BEHAVIORAL of G_GENERAL_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_14 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_14;

architecture SYN_BEHAVIORAL of G_GENERAL_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_340;

architecture SYN_BEHAVIORAL of FA_340 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n3, n_1080 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   MY_CLK_r_REG17_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n3, QN => 
                           n_1080);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3, n7, n_1082 : std_logic;

begin
   
   U7 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   MY_CLK_r_REG80_S2 : DFF_X1 port map( D => n7, CK => clk, Q => n3, QN => 
                           n_1082);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n7, n_1085 : std_logic;

begin
   
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   MY_CLK_r_REG182_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n_1085, QN =>
                           n7);
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n3, n_1087 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   MY_CLK_r_REG183_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n3, QN => 
                           n_1087);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n3, n_1091 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   MY_CLK_r_REG121_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n3, QN => 
                           n_1091);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n7, n_1093 : std_logic;

begin
   
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   MY_CLK_r_REG122_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n_1093, QN =>
                           n7);
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n3, n_1096 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   MY_CLK_r_REG83_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n3, QN => 
                           n_1096);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n_1098 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U7 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   MY_CLK_r_REG82_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n_1098, QN => 
                           n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n_1100 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n8, Z => S);
   MY_CLK_r_REG90_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n_1100, QN => 
                           n8);
   U2 : XNOR2_X1 port map( A => n2, B => n9, ZN => n4);
   U3 : INV_X1 port map( A => B, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2, n4, n3, n7, n_1102 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   MY_CLK_r_REG91_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n3, QN => 
                           n_1102);
   U3 : XNOR2_X1 port map( A => n2, B => n7, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n7, n_1104 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   MY_CLK_r_REG96_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n_1104, QN => 
                           n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n3, n_1106 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   MY_CLK_r_REG97_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n3, QN => 
                           n_1106);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3, n7, n_1108 : std_logic;

begin
   
   U7 : XOR2_X1 port map( A => Ci, B => n3, Z => S);
   MY_CLK_r_REG112_S2 : DFF_X1 port map( D => n7, CK => clk, Q => n3, QN => 
                           n_1108);
   U1 : XOR2_X1 port map( A => A, B => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n1, n2 : std_logic;

begin
   S <= S_port;
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_port);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n3, n_1111 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   MY_CLK_r_REG113_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n3, QN => 
                           n_1111);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_9 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_9;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_9 is

   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X2 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_17 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_17;

architecture SYN_STRUCTURAL of RCA_generic_N2_17 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102704, n_1115 : std_logic;

begin
   
   net102704 <= '0';
   FAI_1 : FA_34 port map( A => A(0), B => B(0), Ci => net102704, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_33 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1115, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_18 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_18;

architecture SYN_STRUCTURAL of RCA_generic_N2_18 is

   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102705, n_1118 : std_logic;

begin
   
   net102705 <= '0';
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => net102705, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1118, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_10 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_10;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_11 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_11;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_12 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_12;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_23 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_23;

architecture SYN_STRUCTURAL of RCA_generic_N2_23 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102706, n_1121 : std_logic;

begin
   
   net102706 <= '0';
   FAI_1 : FA_46 port map( A => A(0), B => B(0), Ci => net102706, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_45 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1121, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_24 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_24;

architecture SYN_STRUCTURAL of RCA_generic_N2_24 is

   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102707, n_1124 : std_logic;

begin
   
   net102707 <= '0';
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => net102707, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1124, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_25 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_25;

architecture SYN_STRUCTURAL of RCA_generic_N2_25 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102701, n_1127 : std_logic;

begin
   
   net102701 <= '0';
   FAI_1 : FA_50 port map( A => A(0), B => B(0), Ci => net102701, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_49 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1127);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_26 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_26;

architecture SYN_STRUCTURAL of RCA_generic_N2_26 is

   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102698, n_1130 : std_logic;

begin
   
   net102698 <= '0';
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => net102698, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1130);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_14 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_14;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_27 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_27;

architecture SYN_STRUCTURAL of RCA_generic_N2_27 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102708, n_1133 : std_logic;

begin
   
   net102708 <= '0';
   FAI_1 : FA_54 port map( A => A(0), B => B(0), Ci => net102708, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_53 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1133);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_28 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_28;

architecture SYN_STRUCTURAL of RCA_generic_N2_28 is

   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102709, n_1136 : std_logic;

begin
   
   net102709 <= '0';
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => net102709, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1136);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_30 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_30;

architecture SYN_STRUCTURAL of RCA_generic_N2_30 is

   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102702, n_1139 : std_logic;

begin
   
   net102702 <= '0';
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => net102702, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1139);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_31 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_31;

architecture SYN_STRUCTURAL of RCA_generic_N2_31 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102703, n_1142 : std_logic;

begin
   
   net102703 <= '0';
   FAI_1 : FA_62 port map( A => A(0), B => B(0), Ci => net102703, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_61 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1142);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_32 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic);

end RCA_generic_N2_32;

architecture SYN_STRUCTURAL of RCA_generic_N2_32 is

   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102711, n_1145 : std_logic;

begin
   
   net102711 <= '0';
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => net102711, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1145);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_33 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_33;

architecture SYN_STRUCTURAL of RCA_generic_N2_33 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102712, n_1148 : std_logic;

begin
   
   net102712 <= '0';
   FAI_1 : FA_66 port map( A => A(0), B => B(0), Ci => net102712, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_65 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1148, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_34 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_34;

architecture SYN_STRUCTURAL of RCA_generic_N2_34 is

   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102713, n_1151 : std_logic;

begin
   
   net102713 <= '0';
   FAI_1 : FA_68 port map( A => A(0), B => B(0), Ci => net102713, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_67 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1151, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_35 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_35;

architecture SYN_STRUCTURAL of RCA_generic_N2_35 is

   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102714, n_1154 : std_logic;

begin
   
   net102714 <= '0';
   FAI_1 : FA_70 port map( A => A(0), B => B(0), Ci => net102714, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_69 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1154, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_36 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_36;

architecture SYN_STRUCTURAL of RCA_generic_N2_36 is

   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102715, n_1157 : std_logic;

begin
   
   net102715 <= '0';
   FAI_1 : FA_72 port map( A => A(0), B => B(0), Ci => net102715, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_71 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1157, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_37 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_37;

architecture SYN_STRUCTURAL of RCA_generic_N2_37 is

   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102716, n_1160 : std_logic;

begin
   
   net102716 <= '0';
   FAI_1 : FA_74 port map( A => A(0), B => B(0), Ci => net102716, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_73 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1160, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_38 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_38;

architecture SYN_STRUCTURAL of RCA_generic_N2_38 is

   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102717, n_1163 : std_logic;

begin
   
   net102717 <= '0';
   FAI_1 : FA_76 port map( A => A(0), B => B(0), Ci => net102717, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_75 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1163, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_39 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_39;

architecture SYN_STRUCTURAL of RCA_generic_N2_39 is

   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102718, n_1166 : std_logic;

begin
   
   net102718 <= '0';
   FAI_1 : FA_78 port map( A => A(0), B => B(0), Ci => net102718, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_77 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1166, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_40 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_40;

architecture SYN_STRUCTURAL of RCA_generic_N2_40 is

   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102719, n_1169 : std_logic;

begin
   
   net102719 <= '0';
   FAI_1 : FA_80 port map( A => A(0), B => B(0), Ci => net102719, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_79 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1169, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N2_21 is

   port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (1 downto 0));

end MUX21_GENERIC_N2_21;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N2_21 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_41 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_41;

architecture SYN_STRUCTURAL of RCA_generic_N2_41 is

   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102720, n_1172 : std_logic;

begin
   
   net102720 <= '0';
   FAI_1 : FA_82 port map( A => A(0), B => B(0), Ci => net102720, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_81 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1172, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N2_42 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
         std_logic);

end RCA_generic_N2_42;

architecture SYN_STRUCTURAL of RCA_generic_N2_42 is

   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_1_port, net102721, n_1175 : std_logic;

begin
   
   net102721 <= '0';
   FAI_1 : FA_84 port map( A => A(0), B => B(0), Ci => net102721, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_83 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => n_1175, clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_9 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_9;

architecture SYN_STRUCTURAL of carry_select_N2_9 is

   component MUX21_GENERIC_N2_9
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_17
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component RCA_generic_N2_18
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n3, n4, n_1176, n_1177, n_1178, n_1179 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG224_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n4, QN => 
                           n_1176);
   MY_CLK_r_REG215_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n3, QN => 
                           n_1177);
   ADDER0 : RCA_generic_N2_18 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1178, clk => clk);
   ADDER1 : RCA_generic_N2_17 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1179, clk => clk);
   MUX : MUX21_GENERIC_N2_9 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_10 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_10;

architecture SYN_STRUCTURAL of carry_select_N2_10 is

   component MUX21_GENERIC_N2_10
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_19
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N2_20
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n2, n_1180, n_1181, n_1182 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG217_S2 : DFF_X1 port map( D => A(1), CK => clk, Q => n2, QN => 
                           n_1180);
   ADDER0 : RCA_generic_N2_20 port map( A(1) => n2, A(0) => A(0), B(1) => B(1),
                           B(0) => B(0), Ci => X_Logic0_port, S(1) => S0_1_port
                           , S(0) => S0_0_port, Co => n_1181);
   ADDER1 : RCA_generic_N2_19 port map( A(1) => n2, A(0) => A(0), B(1) => B(1),
                           B(0) => B(0), Ci => X_Logic1_port, S(1) => S1_1_port
                           , S(0) => S1_0_port, Co => n_1182);
   MUX : MUX21_GENERIC_N2_10 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_11 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_11;

architecture SYN_STRUCTURAL of carry_select_N2_11 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX21_GENERIC_N2_11
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_21
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N2_22
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n5, n6, n7, n8, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG199_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n7, QN => 
                           n_1183);
   MY_CLK_r_REG197_S2 : DFF_X1 port map( D => B(1), CK => clk, Q => n6, QN => 
                           n_1184);
   MY_CLK_r_REG200_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n5, QN => 
                           n_1185);
   ADDER0 : RCA_generic_N2_22 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1186);
   ADDER1 : RCA_generic_N2_21 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1187);
   MUX : MUX21_GENERIC_N2_11 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));
   MY_CLK_r_REG210_S2 : DFF_X1 port map( D => A(1), CK => clk, Q => n8, QN => 
                           n_1188);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_12 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_12;

architecture SYN_STRUCTURAL of carry_select_N2_12 is

   component MUX21_GENERIC_N2_12
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_23
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component RCA_generic_N2_24
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n3, n4, n_1189, n_1190, n_1191, n_1192 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG184_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n4, QN => 
                           n_1189);
   MY_CLK_r_REG188_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n3, QN => 
                           n_1190);
   ADDER0 : RCA_generic_N2_24 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1191, clk => clk);
   ADDER1 : RCA_generic_N2_23 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1192, clk => clk);
   MUX : MUX21_GENERIC_N2_12 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_13 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_13;

architecture SYN_STRUCTURAL of carry_select_N2_13 is

   component MUX21_GENERIC_N2_13
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_25
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N2_26
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n5, n6, n7, n8, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG187_S2 : DFF_X1 port map( D => A(1), CK => clk, Q => n8, QN => 
                           n_1193);
   MY_CLK_r_REG168_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n7, QN => 
                           n_1194);
   MY_CLK_r_REG165_S2 : DFF_X1 port map( D => B(1), CK => clk, Q => n6, QN => 
                           n_1195);
   MY_CLK_r_REG171_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n5, QN => 
                           n_1196);
   ADDER0 : RCA_generic_N2_26 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1197);
   ADDER1 : RCA_generic_N2_25 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1198);
   MUX : MUX21_GENERIC_N2_13 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_14 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_14;

architecture SYN_STRUCTURAL of carry_select_N2_14 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX21_GENERIC_N2_14
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_27
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N2_28
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n5, n6, n7, n8, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG154_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n7, QN => 
                           n_1199);
   MY_CLK_r_REG152_S2 : DFF_X1 port map( D => B(1), CK => clk, Q => n6, QN => 
                           n_1200);
   MY_CLK_r_REG156_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n5, QN => 
                           n_1201);
   ADDER0 : RCA_generic_N2_28 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1202);
   ADDER1 : RCA_generic_N2_27 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1203);
   MUX : MUX21_GENERIC_N2_14 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));
   MY_CLK_r_REG170_S2 : DFF_X1 port map( D => A(1), CK => clk, Q => n8, QN => 
                           n_1204);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_15 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_15;

architecture SYN_STRUCTURAL of carry_select_N2_15 is

   component MUX21_GENERIC_N2_15
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_29
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N2_30
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n5, n6, n7, n8, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG155_S2 : DFF_X1 port map( D => A(1), CK => clk, Q => n8, QN => 
                           n_1205);
   MY_CLK_r_REG142_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n7, QN => 
                           n_1206);
   MY_CLK_r_REG140_S2 : DFF_X1 port map( D => B(1), CK => clk, Q => n6, QN => 
                           n_1207);
   MY_CLK_r_REG128_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n5, QN => 
                           n_1208);
   ADDER0 : RCA_generic_N2_30 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1209);
   ADDER1 : RCA_generic_N2_29 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1210);
   MUX : MUX21_GENERIC_N2_15 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_16 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_16;

architecture SYN_STRUCTURAL of carry_select_N2_16 is

   component MUX21_GENERIC_N2_16
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_31
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N2_32
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n5, n6, n7, n8, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216
      : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG131_S2 : DFF_X1 port map( D => A(1), CK => clk, Q => n8, QN => 
                           n_1211);
   MY_CLK_r_REG134_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n7, QN => 
                           n_1212);
   MY_CLK_r_REG133_S2 : DFF_X1 port map( D => B(1), CK => clk, Q => n6, QN => 
                           n_1213);
   MY_CLK_r_REG120_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n5, QN => 
                           n_1214);
   ADDER0 : RCA_generic_N2_32 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1215);
   ADDER1 : RCA_generic_N2_31 port map( A(1) => n8, A(0) => n7, B(1) => n6, 
                           B(0) => n5, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1216);
   MUX : MUX21_GENERIC_N2_16 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_17 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_17;

architecture SYN_STRUCTURAL of carry_select_N2_17 is

   component MUX21_GENERIC_N2_17
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_33
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component RCA_generic_N2_34
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n3, n4, n_1217, n_1218, n_1219, n_1220 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG123_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n4, QN => 
                           n_1217);
   MY_CLK_r_REG104_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n3, QN => 
                           n_1218);
   ADDER0 : RCA_generic_N2_34 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1219, clk => clk);
   ADDER1 : RCA_generic_N2_33 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1220, clk => clk);
   MUX : MUX21_GENERIC_N2_17 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_18 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_18;

architecture SYN_STRUCTURAL of carry_select_N2_18 is

   component MUX21_GENERIC_N2_18
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_35
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component RCA_generic_N2_36
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n3, n4, n_1221, n_1222, n_1223, n_1224 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG87_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n4, QN => 
                           n_1221);
   MY_CLK_r_REG89_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n3, QN => 
                           n_1222);
   ADDER0 : RCA_generic_N2_36 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1223, clk => clk);
   ADDER1 : RCA_generic_N2_35 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1224, clk => clk);
   MUX : MUX21_GENERIC_N2_18 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_19 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_19;

architecture SYN_STRUCTURAL of carry_select_N2_19 is

   component MUX21_GENERIC_N2_19
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_37
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component RCA_generic_N2_38
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n3, n4, n_1225, n_1226, n_1227, n_1228 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG94_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n4, QN => 
                           n_1225);
   MY_CLK_r_REG95_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n3, QN => 
                           n_1226);
   ADDER0 : RCA_generic_N2_38 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1227, clk => clk);
   ADDER1 : RCA_generic_N2_37 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1228, clk => clk);
   MUX : MUX21_GENERIC_N2_19 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_20 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_20;

architecture SYN_STRUCTURAL of carry_select_N2_20 is

   component MUX21_GENERIC_N2_20
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_39
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component RCA_generic_N2_40
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n3, n4, n_1229, n_1230, n_1231, n_1232 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG102_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n4, QN => 
                           n_1229);
   MY_CLK_r_REG116_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n3, QN => 
                           n_1230);
   ADDER0 : RCA_generic_N2_40 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1231, clk => clk);
   ADDER1 : RCA_generic_N2_39 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1232, clk => clk);
   MUX : MUX21_GENERIC_N2_20 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N2_21 is

   port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end carry_select_N2_21;

architecture SYN_STRUCTURAL of carry_select_N2_21 is

   component MUX21_GENERIC_N2_21
      port( A, B : in std_logic_vector (1 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (1 downto 0));
   end component;
   
   component RCA_generic_N2_41
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component RCA_generic_N2_42
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_1_port, S0_0_port, S1_1_port, 
      S1_0_port, n3, n4, n_1233, n_1234, n_1235, n_1236 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG266_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n4, QN => 
                           n_1233);
   MY_CLK_r_REG279_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n3, QN => 
                           n_1234);
   ADDER0 : RCA_generic_N2_42 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic0_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1235, clk => clk);
   ADDER1 : RCA_generic_N2_41 port map( A(1) => A(1), A(0) => n4, B(1) => B(1),
                           B(0) => n3, Ci => X_Logic1_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1236, clk => clk);
   MUX : MUX21_GENERIC_N2_21 port map( A(1) => S1_1_port, A(0) => S1_0_port, 
                           B(1) => S0_1_port, B(0) => S0_0_port, SEL => Ci, 
                           Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_10 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_10;

architecture SYN_BEHAVIORAL of G_GENERAL_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_11 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_11;

architecture SYN_BEHAVIORAL of G_GENERAL_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_12 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_12;

architecture SYN_BEHAVIORAL of G_GENERAL_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_17 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_17;

architecture SYN_BEHAVIORAL of G_GENERAL_17 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => G_k_1j, A2 => PG_ik(0), ZN => n2);
   U1 : OR2_X1 port map( A1 => PG_ik(1), A2 => n2, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_21 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_21;

architecture SYN_BEHAVIORAL of G_GENERAL_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_14 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_14;

architecture SYN_BEHAVIORAL of PG_GENERAL_14 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => PG_ik(1), A2 => PG_ik(0), ZN => n2);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => PG_ij(1));
   U4 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : NOR2_X1 port map( A1 => PG_ik(1), A2 => PG_k_1j(1), ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_15 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_15;

architecture SYN_BEHAVIORAL of PG_GENERAL_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_16 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_16;

architecture SYN_BEHAVIORAL of PG_GENERAL_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_17 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_17;

architecture SYN_BEHAVIORAL of PG_GENERAL_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => PG_ik(1), A2 => n2, ZN => PG_ij(1));
   U2 : AND2_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(0), ZN => n2);
   U3 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_19 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_19;

architecture SYN_BEHAVIORAL of PG_GENERAL_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_20 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_20;

architecture SYN_BEHAVIORAL of PG_GENERAL_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_25 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic;  clk : in std_logic);

end G_GENERAL_25;

architecture SYN_BEHAVIORAL of G_GENERAL_25 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n_1237 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   MY_CLK_r_REG344_S2 : DFF_X1 port map( D => n1, CK => clk, Q => n_1237, QN =>
                           G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_27 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_27;

architecture SYN_BEHAVIORAL of PG_GENERAL_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_29 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_29;

architecture SYN_BEHAVIORAL of PG_GENERAL_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U4 : INV_X1 port map( A => n2, ZN => PG_ij(1));
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_31 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_31;

architecture SYN_BEHAVIORAL of PG_GENERAL_31 is

   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n_1238, n_1239 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => PG_k_1j(1), A2 => n4, ZN => n2);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => n4, ZN => PG_ij(0));
   MY_CLK_r_REG114_S2 : DFF_X1 port map( D => PG_ik(1), CK => clk, Q => n5, QN 
                           => n_1238);
   MY_CLK_r_REG115_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n4, QN 
                           => n_1239);
   U1 : OR2_X2 port map( A1 => n2, A2 => n5, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_32 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_32;

architecture SYN_BEHAVIORAL of PG_GENERAL_32 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n5, n_1240, n_1241 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => n4, ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => n4, A => n5, ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   MY_CLK_r_REG277_S2 : DFF_X1 port map( D => PG_ik(1), CK => clk, Q => n5, QN 
                           => n_1240);
   MY_CLK_r_REG278_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n4, QN 
                           => n_1241);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_29 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_29;

architecture SYN_BEHAVIORAL of G_GENERAL_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_41 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_41;

architecture SYN_BEHAVIORAL of PG_GENERAL_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_42 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_42;

architecture SYN_BEHAVIORAL of PG_GENERAL_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_43 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_43;

architecture SYN_BEHAVIORAL of PG_GENERAL_43 is

   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n6, n9, n10, n11, n_1242 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n6, A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : OAI21_X1 port map( B1 => n3, B2 => n11, A => n9, ZN => PG_ij(1));
   U3 : INV_X1 port map( A => PG_k_1j(1), ZN => n3);
   MY_CLK_r_REG106_S2 : DFF_X1 port map( D => PG_ik(1), CK => clk, Q => n_1242,
                           QN => n9);
   MY_CLK_r_REG105_S2 : DFFS_X1 port map( D => PG_ik(0), CK => clk, SN => n10, 
                           Q => n6, QN => n11);
   n10 <= '1';

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_44 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_44;

architecture SYN_BEHAVIORAL of PG_GENERAL_44 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n5, n_1243, n_1244 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => n4, ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => n4, A => n5, ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   MY_CLK_r_REG93_S2 : DFF_X1 port map( D => PG_ik(1), CK => clk, Q => n5, QN 
                           => n_1243);
   MY_CLK_r_REG92_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n4, QN 
                           => n_1244);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_31 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic;  clk : in std_logic);

end G_GENERAL_31;

architecture SYN_BEHAVIORAL of G_GENERAL_31 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n_1245 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   MY_CLK_r_REG451_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n_1245, QN =>
                           G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_59 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_59;

architecture SYN_BEHAVIORAL of PG_GENERAL_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => PG_ik(1), ZN => n3);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => PG_ij(1));
   U4 : NAND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_60 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_60;

architecture SYN_BEHAVIORAL of PG_GENERAL_60 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n6, n7, n_1246, n_1247, n_1248 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n6, A2 => n7, ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   MY_CLK_r_REG195_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n7, QN 
                           => n_1246);
   MY_CLK_r_REG198_S2 : DFF_X1 port map( D => PG_k_1j(0), CK => clk, Q => n6, 
                           QN => n_1247);
   MY_CLK_r_REG196_S2 : DFF_X1 port map( D => n1, CK => clk, Q => n_1248, QN =>
                           PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_61 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_61;

architecture SYN_BEHAVIORAL of PG_GENERAL_61 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n8, n12, n13, n14, n_1249, n_1250, n_1251 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n6, A2 => n8, ZN => PG_ij(0));
   MY_CLK_r_REG186_S2 : DFF_X1 port map( D => PG_k_1j(0), CK => clk, Q => n6, 
                           QN => n_1249);
   MY_CLK_r_REG185_S2 : DFF_X1 port map( D => PG_k_1j(1), CK => clk, Q => 
                           n_1250, QN => n12);
   MY_CLK_r_REG180_S2 : DFF_X1 port map( D => PG_ik(1), CK => clk, Q => n_1251,
                           QN => n14);
   U2 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n14, ZN => PG_ij(1));
   MY_CLK_r_REG181_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n8, QN 
                           => n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_62 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_62;

architecture SYN_BEHAVIORAL of PG_GENERAL_62 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n6, n7, n_1252, n_1253, n_1254 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : AND2_X1 port map( A1 => n7, A2 => n6, ZN => PG_ij(0));
   MY_CLK_r_REG169_S2 : DFF_X1 port map( D => PG_k_1j(0), CK => clk, Q => n6, 
                           QN => n_1252);
   MY_CLK_r_REG166_S2 : DFF_X1 port map( D => n1, CK => clk, Q => n_1253, QN =>
                           PG_ij(1));
   MY_CLK_r_REG167_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n7, QN 
                           => n_1254);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_63 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_63;

architecture SYN_BEHAVIORAL of PG_GENERAL_63 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n6, n7, n_1255, n_1256, n_1257 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n6, A2 => n7, ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   MY_CLK_r_REG153_S2 : DFF_X1 port map( D => PG_k_1j(0), CK => clk, Q => n6, 
                           QN => n_1255);
   MY_CLK_r_REG150_S2 : DFF_X1 port map( D => n1, CK => clk, Q => n_1256, QN =>
                           PG_ij(1));
   MY_CLK_r_REG151_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n7, QN 
                           => n_1257);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_64 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_64;

architecture SYN_BEHAVIORAL of PG_GENERAL_64 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n6, n7, n_1258, n_1259, n_1260 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n7, A2 => n6, ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   MY_CLK_r_REG141_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n7, QN 
                           => n_1258);
   MY_CLK_r_REG130_S2 : DFF_X1 port map( D => PG_k_1j(0), CK => clk, Q => n6, 
                           QN => n_1259);
   MY_CLK_r_REG129_S2 : DFF_X1 port map( D => n1, CK => clk, Q => n_1260, QN =>
                           PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_65 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_65;

architecture SYN_BEHAVIORAL of PG_GENERAL_65 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n_1261, n_1262 : std_logic;

begin
   
   U4 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => n5, ZN => PG_ij(0));
   U1 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   MY_CLK_r_REG132_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n5, QN 
                           => n_1261);
   MY_CLK_r_REG119_S2 : DFF_X1 port map( D => n1, CK => clk, Q => n_1262, QN =>
                           PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_66 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_66;

architecture SYN_BEHAVIORAL of PG_GENERAL_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => PG_ik(1), ZN => n6);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => PG_ij(1));
   U4 : NAND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_67 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_67;

architecture SYN_BEHAVIORAL of PG_GENERAL_67 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n7, n8, n9, n_1263, n_1264, n_1265 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : OAI21_X1 port map( B1 => n9, B2 => n8, A => n7, ZN => PG_ij(1));
   U3 : INV_X1 port map( A => PG_ik(0), ZN => n3);
   U4 : INV_X1 port map( A => PG_k_1j(1), ZN => n4);
   U5 : INV_X1 port map( A => PG_ik(1), ZN => n5);
   MY_CLK_r_REG86_S2 : DFF_X1 port map( D => n3, CK => clk, Q => n9, QN => 
                           n_1263);
   MY_CLK_r_REG88_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n8, QN => 
                           n_1264);
   MY_CLK_r_REG84_S2 : DFF_X1 port map( D => n5, CK => clk, Q => n7, QN => 
                           n_1265);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_70 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_70;

architecture SYN_BEHAVIORAL of PG_GENERAL_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_72 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_72;

architecture SYN_BEHAVIORAL of PG_GENERAL_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_74 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_74;

architecture SYN_BEHAVIORAL of PG_GENERAL_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_77 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_77;

architecture SYN_BEHAVIORAL of PG_GENERAL_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_0 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_0;

architecture SYN_BEHAVIORAL of PG_GENERAL_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_0 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_0;

architecture SYN_BEHAVIORAL of G_GENERAL_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => G_k_1j, A2 => PG_ik(0), ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_19 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
         std_logic);

end PG_NET_19;

architecture SYN_BEHAVIORAL of PG_NET_19 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n_1267 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n4, A2 => n1, ZN => G_OUT);
   MY_CLK_r_REG216_S2 : DFF_X1 port map( D => n2, CK => clk, Q => n4, QN => 
                           n_1267);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_25 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_25;

architecture SYN_BEHAVIORAL of PG_NET_25 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net29650, net29651 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => net29650);
   U3 : INV_X1 port map( A => B, ZN => net29651);
   U4 : NOR2_X1 port map( A1 => net29650, A2 => net29651, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_26 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_26;

architecture SYN_BEHAVIORAL of PG_NET_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_27 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_27;

architecture SYN_BEHAVIORAL of PG_NET_27 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_29 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_29;

architecture SYN_BEHAVIORAL of PG_NET_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_31 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_31;

architecture SYN_BEHAVIORAL of PG_NET_31 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net29662, net29663 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => net29662);
   U3 : INV_X1 port map( A => B, ZN => net29663);
   U4 : NOR2_X1 port map( A1 => net29662, A2 => net29663, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_32 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
         std_logic);

end PG_NET_32;

architecture SYN_BEHAVIORAL of PG_NET_32 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n_1268, n_1269 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U3 : XOR2_X1 port map( A => n4, B => n5, Z => P_OUT);
   MY_CLK_r_REG135_S2 : DFF_X1 port map( D => A, CK => clk, Q => n5, QN => 
                           n_1268);
   MY_CLK_r_REG118_S2 : DFF_X1 port map( D => B, CK => clk, Q => n4, QN => 
                           n_1269);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_35 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_35;

architecture SYN_BEHAVIORAL of PG_NET_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_37 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_37;

architecture SYN_BEHAVIORAL of PG_NET_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U3 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_38 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_38;

architecture SYN_BEHAVIORAL of PG_NET_38 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : INV_X1 port map( A => B, ZN => n1);
   U3 : XNOR2_X1 port map( A => A, B => n1, ZN => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_42 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_42;

architecture SYN_BEHAVIORAL of PG_NET_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_44 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_44;

architecture SYN_BEHAVIORAL of PG_NET_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_45 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_45;

architecture SYN_BEHAVIORAL of PG_NET_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_49 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_49;

architecture SYN_BEHAVIORAL of PG_NET_49 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_50 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_50;

architecture SYN_BEHAVIORAL of PG_NET_50 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_52 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_52;

architecture SYN_BEHAVIORAL of PG_NET_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_53 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_53;

architecture SYN_BEHAVIORAL of PG_NET_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_54 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_54;

architecture SYN_BEHAVIORAL of PG_NET_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_58 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
         std_logic);

end PG_NET_58;

architecture SYN_BEHAVIORAL of PG_NET_58 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n_1270 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => n2, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => n2, B => A, Z => P_OUT);
   MY_CLK_r_REG436_S1 : DFF_X1 port map( D => B, CK => clk, Q => n2, QN => 
                           n_1270);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_59 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
         std_logic);

end PG_NET_59;

architecture SYN_BEHAVIORAL of PG_NET_59 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6, n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n5, B => n6, Z => P_OUT);
   U4 : NOR2_X1 port map( A1 => n8, A2 => n9, ZN => G_OUT);
   MY_CLK_r_REG437_S1 : DFF_X1 port map( D => A, CK => clk, Q => n6, QN => n8);
   MY_CLK_r_REG447_S1 : DFF_X1 port map( D => B, CK => clk, Q => n5, QN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_60 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
         std_logic);

end PG_NET_60;

architecture SYN_BEHAVIORAL of PG_NET_60 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n5, n6, n8, n9 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n5, B => n6, Z => P_OUT);
   U4 : NOR2_X1 port map( A1 => n9, A2 => n8, ZN => G_OUT);
   MY_CLK_r_REG452_S1 : DFF_X1 port map( D => B, CK => clk, Q => n5, QN => n8);
   MY_CLK_r_REG448_S1 : DFF_X1 port map( D => A, CK => clk, Q => n6, QN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_62 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_62;

architecture SYN_BEHAVIORAL of PG_NET_62 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_63 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_63;

architecture SYN_BEHAVIORAL of PG_NET_63 is

begin
   P_OUT <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_0 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_0;

architecture SYN_BEHAVIORAL of PG_NET_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK2_NBLOCKS32 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic_vector 
         (31 downto 0);  S : out std_logic_vector (63 downto 0);  clk : in 
         std_logic);

end SUM_GENERATOR_NBIT_PER_BLOCK2_NBLOCKS32;

architecture SYN_STRUCTURAL of SUM_GENERATOR_NBIT_PER_BLOCK2_NBLOCKS32 is

   component carry_select_N2_9
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_10
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_11
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_12
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_13
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_14
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_15
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_16
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_17
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_18
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_19
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_20
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N2_21
      port( A, B : in std_logic_vector (1 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;

begin
   
   CS_11 : carry_select_N2_21 port map( A(1) => A(23), A(0) => A(22), B(1) => 
                           B(23), B(0) => B(22), Ci => Ci(11), S(1) => S(23), 
                           S(0) => S(22), clk => clk);
   CS_12 : carry_select_N2_20 port map( A(1) => A(25), A(0) => A(24), B(1) => 
                           B(25), B(0) => B(24), Ci => Ci(12), S(1) => S(25), 
                           S(0) => S(24), clk => clk);
   CS_13 : carry_select_N2_19 port map( A(1) => A(27), A(0) => A(26), B(1) => 
                           B(27), B(0) => B(26), Ci => Ci(13), S(1) => S(27), 
                           S(0) => S(26), clk => clk);
   CS_14 : carry_select_N2_18 port map( A(1) => A(29), A(0) => A(28), B(1) => 
                           B(29), B(0) => B(28), Ci => Ci(14), S(1) => S(29), 
                           S(0) => S(28), clk => clk);
   CS_15 : carry_select_N2_17 port map( A(1) => A(31), A(0) => A(30), B(1) => 
                           B(31), B(0) => B(30), Ci => Ci(15), S(1) => S(31), 
                           S(0) => S(30), clk => clk);
   CS_16 : carry_select_N2_16 port map( A(1) => A(33), A(0) => A(32), B(1) => 
                           B(33), B(0) => B(32), Ci => Ci(16), S(1) => S(33), 
                           S(0) => S(32), clk => clk);
   CS_17 : carry_select_N2_15 port map( A(1) => A(35), A(0) => A(34), B(1) => 
                           B(35), B(0) => B(34), Ci => Ci(17), S(1) => S(35), 
                           S(0) => S(34), clk => clk);
   CS_18 : carry_select_N2_14 port map( A(1) => A(37), A(0) => A(36), B(1) => 
                           B(37), B(0) => B(36), Ci => Ci(18), S(1) => S(37), 
                           S(0) => S(36), clk => clk);
   CS_19 : carry_select_N2_13 port map( A(1) => A(39), A(0) => A(38), B(1) => 
                           B(39), B(0) => B(38), Ci => Ci(19), S(1) => S(39), 
                           S(0) => S(38), clk => clk);
   CS_20 : carry_select_N2_12 port map( A(1) => A(41), A(0) => A(40), B(1) => 
                           B(41), B(0) => B(40), Ci => Ci(20), S(1) => S(41), 
                           S(0) => S(40), clk => clk);
   CS_21 : carry_select_N2_11 port map( A(1) => A(43), A(0) => A(42), B(1) => 
                           B(43), B(0) => B(42), Ci => Ci(21), S(1) => S(43), 
                           S(0) => S(42), clk => clk);
   CS_22 : carry_select_N2_10 port map( A(1) => A(45), A(0) => A(44), B(1) => 
                           B(45), B(0) => B(44), Ci => Ci(22), S(1) => S(45), 
                           S(0) => S(44), clk => clk);
   CS_23 : carry_select_N2_9 port map( A(1) => A(47), A(0) => A(46), B(1) => 
                           B(47), B(0) => B(46), Ci => Ci(23), S(1) => S(47), 
                           S(0) => S(46), clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK2 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (32 downto 0);  clk : in std_logic);

end CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK2;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK2 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component G_GENERAL_10
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_11
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_12
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_13
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_14
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_15
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_16
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_17
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_18
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_19
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_20
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_21
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_22
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_14
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_15
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_16
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_17
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_18
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_19
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_20
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_25
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic;  clk : in std_logic);
   end component;
   
   component PG_GENERAL_26
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_27
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_28
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_29
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_30
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_31
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_32
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_33
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_29
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_40
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_41
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_42
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_43
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_44
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_45
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_46
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_47
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_48
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_49
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_31
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic;  clk : in std_logic);
   end component;
   
   component PG_GENERAL_59
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_60
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_61
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_62
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_63
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_64
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_65
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_66
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_67
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_68
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_69
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_70
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_71
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_72
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_73
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_74
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_75
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_76
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_77
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_78
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_79
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_0
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_0
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_NET_19
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component PG_NET_20
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_21
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_22
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_23
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_24
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_25
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_26
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_27
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_28
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_29
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_30
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_31
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_32
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component PG_NET_33
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_34
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_35
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_36
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_37
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_38
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_39
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_40
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_41
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_42
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_43
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_44
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_45
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_46
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_47
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_48
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_49
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_50
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_51
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_52
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_53
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_54
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_55
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_56
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_57
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_58
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component PG_NET_59
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component PG_NET_60
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component PG_NET_61
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_62
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_63
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_0
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   signal Co_22_port, Co_21_port, Co_20_port, Co_19_port, Co_18_port, 
      Co_17_port, n16, Co_15_port, Co_14_port, Co_13_port, Co_12_port, 
      Co_11_port, n17, n25, n26, n27, lev_i_out_4_46_1_port, 
      lev_i_out_4_46_0_port, lev_i_out_4_44_1_port, lev_i_out_4_44_0_port, 
      lev_i_out_4_42_1_port, lev_i_out_4_42_0_port, lev_i_out_4_32_1_port, 
      lev_i_out_4_32_0_port, lev_i_out_4_30_1_port, lev_i_out_4_30_0_port, 
      lev_i_out_4_28_1_port, lev_i_out_4_28_0_port, lev_i_out_4_26_1_port, 
      lev_i_out_4_26_0_port, lev_i_out_3_46_1_port, lev_i_out_3_46_0_port, 
      lev_i_out_3_40_0_port, lev_i_out_3_38_1_port, lev_i_out_3_38_0_port, 
      lev_i_out_3_32_1_port, lev_i_out_3_32_0_port, lev_i_out_3_30_1_port, 
      lev_i_out_3_30_0_port, lev_i_out_3_24_0_port, lev_i_out_3_22_1_port, 
      lev_i_out_3_22_0_port, lev_i_out_3_16_1_port, lev_i_out_3_16_0_port, 
      lev_i_out_2_44_1_port, lev_i_out_2_44_0_port, lev_i_out_2_40_1_port, 
      lev_i_out_2_40_0_port, lev_i_out_2_36_1_port, lev_i_out_2_36_0_port, 
      lev_i_out_2_32_1_port, lev_i_out_2_32_0_port, lev_i_out_2_28_1_port, 
      lev_i_out_2_28_0_port, lev_i_out_2_24_1_port, lev_i_out_2_24_0_port, 
      lev_i_out_2_20_1_port, lev_i_out_2_20_0_port, lev_i_out_2_16_1_port, 
      lev_i_out_2_16_0_port, lev_i_out_2_12_1_port, lev_i_out_2_12_0_port, 
      lev_i_out_2_8_1_port, lev_i_out_2_8_0_port, lev_i_out_1_46_1_port, 
      lev_i_out_1_46_0_port, lev_i_out_1_44_1_port, lev_i_out_1_44_0_port, 
      lev_i_out_1_42_1_port, lev_i_out_1_42_0_port, lev_i_out_1_40_1_port, 
      lev_i_out_1_40_0_port, lev_i_out_1_38_1_port, lev_i_out_1_38_0_port, 
      lev_i_out_1_36_1_port, lev_i_out_1_36_0_port, lev_i_out_1_34_1_port, 
      lev_i_out_1_34_0_port, lev_i_out_1_32_1_port, lev_i_out_1_32_0_port, 
      lev_i_out_1_30_1_port, lev_i_out_1_30_0_port, lev_i_out_1_28_1_port, 
      lev_i_out_1_28_0_port, lev_i_out_1_26_1_port, lev_i_out_1_26_0_port, 
      lev_i_out_1_24_1_port, lev_i_out_1_24_0_port, lev_i_out_1_22_1_port, 
      lev_i_out_1_22_0_port, lev_i_out_1_20_1_port, lev_i_out_1_20_0_port, 
      lev_i_out_1_18_1_port, lev_i_out_1_18_0_port, lev_i_out_1_16_1_port, 
      lev_i_out_1_16_0_port, lev_i_out_1_14_1_port, lev_i_out_1_14_0_port, 
      lev_i_out_1_12_1_port, lev_i_out_1_12_0_port, lev_i_out_1_10_1_port, 
      lev_i_out_1_10_0_port, lev_i_out_1_8_1_port, lev_i_out_1_8_0_port, 
      lev_i_out_1_6_1_port, lev_i_out_1_6_0_port, lev_i_out_1_4_1_port, 
      lev_i_out_1_4_0_port, lev_i_out_0_46_1_port, lev_i_out_0_46_0_port, 
      lev_i_out_0_45_1_port, lev_i_out_0_45_0_port, lev_i_out_0_44_1_port, 
      lev_i_out_0_44_0_port, lev_i_out_0_43_1_port, lev_i_out_0_43_0_port, 
      lev_i_out_0_42_1_port, lev_i_out_0_42_0_port, lev_i_out_0_41_1_port, 
      lev_i_out_0_41_0_port, lev_i_out_0_40_1_port, lev_i_out_0_40_0_port, 
      lev_i_out_0_39_1_port, lev_i_out_0_39_0_port, lev_i_out_0_38_1_port, 
      lev_i_out_0_38_0_port, lev_i_out_0_37_1_port, lev_i_out_0_37_0_port, 
      lev_i_out_0_36_1_port, lev_i_out_0_36_0_port, lev_i_out_0_35_1_port, 
      lev_i_out_0_35_0_port, lev_i_out_0_34_1_port, lev_i_out_0_33_1_port, 
      lev_i_out_0_33_0_port, lev_i_out_0_32_1_port, lev_i_out_0_32_0_port, 
      lev_i_out_0_31_1_port, lev_i_out_0_31_0_port, lev_i_out_0_30_1_port, 
      lev_i_out_0_30_0_port, lev_i_out_0_29_1_port, lev_i_out_0_29_0_port, 
      lev_i_out_0_28_1_port, lev_i_out_0_28_0_port, lev_i_out_0_27_1_port, 
      lev_i_out_0_27_0_port, lev_i_out_0_26_1_port, lev_i_out_0_26_0_port, 
      lev_i_out_0_25_1_port, lev_i_out_0_25_0_port, lev_i_out_0_24_1_port, 
      lev_i_out_0_24_0_port, lev_i_out_0_23_1_port, lev_i_out_0_23_0_port, 
      lev_i_out_0_22_1_port, lev_i_out_0_22_0_port, lev_i_out_0_21_1_port, 
      lev_i_out_0_21_0_port, lev_i_out_0_20_1_port, lev_i_out_0_20_0_port, 
      lev_i_out_0_19_1_port, lev_i_out_0_19_0_port, lev_i_out_0_18_1_port, 
      lev_i_out_0_18_0_port, lev_i_out_0_17_1_port, lev_i_out_0_17_0_port, 
      lev_i_out_0_16_1_port, lev_i_out_0_16_0_port, lev_i_out_0_15_1_port, 
      lev_i_out_0_15_0_port, lev_i_out_0_14_1_port, lev_i_out_0_14_0_port, 
      lev_i_out_0_13_1_port, lev_i_out_0_13_0_port, lev_i_out_0_12_1_port, 
      lev_i_out_0_12_0_port, lev_i_out_0_11_1_port, lev_i_out_0_11_0_port, 
      lev_i_out_0_10_1_port, lev_i_out_0_10_0_port, lev_i_out_0_9_1_port, 
      lev_i_out_0_9_0_port, lev_i_out_0_8_1_port, lev_i_out_0_8_0_port, 
      lev_i_out_0_7_1_port, lev_i_out_0_7_0_port, lev_i_out_0_6_1_port, 
      lev_i_out_0_6_0_port, lev_i_out_0_5_1_port, lev_i_out_0_5_0_port, 
      lev_i_out_0_4_1_port, lev_i_out_0_4_0_port, lev_i_out_0_3_1_port, 
      lev_i_out_0_3_0_port, lev_i_out_0_2_0_port, lev_i_out_0_1_1_port, n19, 
      n20, n21, n22, n23, n28, n30, Co_23_port, n38, net102722, net102723, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471 : 
      std_logic;

begin
   Co <= ( n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, 
      n_1453, Co_23_port, Co_22_port, Co_21_port, Co_20_port, Co_19_port, 
      Co_18_port, Co_17_port, n16, Co_15_port, Co_14_port, Co_13_port, 
      Co_12_port, Co_11_port, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, 
      n_1460, n_1461, n_1462, n_1463, n_1464 );
   
   MY_CLK_r_REG98_S2 : DFF_X1 port map( D => lev_i_out_1_26_1_port, CK => clk, 
                           Q => n23, QN => n_1465);
   MY_CLK_r_REG99_S2 : DFF_X1 port map( D => lev_i_out_1_26_0_port, CK => clk, 
                           Q => n22, QN => n_1466);
   MY_CLK_r_REG300_S2 : DFF_X1 port map( D => lev_i_out_2_20_1_port, CK => clk,
                           Q => n20, QN => n_1467);
   MY_CLK_r_REG301_S2 : DFF_X1 port map( D => lev_i_out_2_20_0_port, CK => clk,
                           Q => n19, QN => n_1468);
   net102722 <= '0';
   net102723 <= '0';
   PG_NETWORK_0_1 : PG_NET_0 port map( A => A(0), B => B(0), G_OUT => 
                           lev_i_out_0_1_1_port, P_OUT => n_1469);
   PG_NETWORK_0_2 : PG_NET_63 port map( A => A(1), B => net102723, G_OUT => 
                           n_1470, P_OUT => lev_i_out_0_2_0_port);
   PG_NETWORK_0_3 : PG_NET_62 port map( A => A(2), B => B(2), G_OUT => 
                           lev_i_out_0_3_1_port, P_OUT => lev_i_out_0_3_0_port)
                           ;
   PG_NETWORK_0_4 : PG_NET_61 port map( A => A(3), B => B(3), G_OUT => 
                           lev_i_out_0_4_1_port, P_OUT => lev_i_out_0_4_0_port)
                           ;
   PG_NETWORK_0_5 : PG_NET_60 port map( A => A(4), B => B(4), G_OUT => 
                           lev_i_out_0_5_1_port, P_OUT => lev_i_out_0_5_0_port,
                           clk => clk);
   PG_NETWORK_0_6 : PG_NET_59 port map( A => A(5), B => B(5), G_OUT => 
                           lev_i_out_0_6_1_port, P_OUT => lev_i_out_0_6_0_port,
                           clk => clk);
   PG_NETWORK_0_7 : PG_NET_58 port map( A => A(6), B => B(6), G_OUT => 
                           lev_i_out_0_7_1_port, P_OUT => lev_i_out_0_7_0_port,
                           clk => clk);
   PG_NETWORK_0_8 : PG_NET_57 port map( A => A(7), B => B(7), G_OUT => 
                           lev_i_out_0_8_1_port, P_OUT => lev_i_out_0_8_0_port)
                           ;
   PG_NETWORK_0_9 : PG_NET_56 port map( A => A(8), B => B(8), G_OUT => 
                           lev_i_out_0_9_1_port, P_OUT => lev_i_out_0_9_0_port)
                           ;
   PG_NETWORK_0_10 : PG_NET_55 port map( A => A(9), B => B(9), G_OUT => 
                           lev_i_out_0_10_1_port, P_OUT => 
                           lev_i_out_0_10_0_port);
   PG_NETWORK_0_11 : PG_NET_54 port map( A => A(10), B => B(10), G_OUT => 
                           lev_i_out_0_11_1_port, P_OUT => 
                           lev_i_out_0_11_0_port);
   PG_NETWORK_0_12 : PG_NET_53 port map( A => A(11), B => B(11), G_OUT => 
                           lev_i_out_0_12_1_port, P_OUT => 
                           lev_i_out_0_12_0_port);
   PG_NETWORK_0_13 : PG_NET_52 port map( A => A(12), B => B(12), G_OUT => 
                           lev_i_out_0_13_1_port, P_OUT => 
                           lev_i_out_0_13_0_port);
   PG_NETWORK_0_14 : PG_NET_51 port map( A => A(13), B => B(13), G_OUT => 
                           lev_i_out_0_14_1_port, P_OUT => 
                           lev_i_out_0_14_0_port);
   PG_NETWORK_0_15 : PG_NET_50 port map( A => A(14), B => B(14), G_OUT => 
                           lev_i_out_0_15_1_port, P_OUT => 
                           lev_i_out_0_15_0_port);
   PG_NETWORK_0_16 : PG_NET_49 port map( A => A(15), B => B(15), G_OUT => 
                           lev_i_out_0_16_1_port, P_OUT => 
                           lev_i_out_0_16_0_port);
   PG_NETWORK_0_17 : PG_NET_48 port map( A => A(16), B => B(16), G_OUT => 
                           lev_i_out_0_17_1_port, P_OUT => 
                           lev_i_out_0_17_0_port);
   PG_NETWORK_0_18 : PG_NET_47 port map( A => A(17), B => B(17), G_OUT => 
                           lev_i_out_0_18_1_port, P_OUT => 
                           lev_i_out_0_18_0_port);
   PG_NETWORK_0_19 : PG_NET_46 port map( A => A(18), B => B(18), G_OUT => 
                           lev_i_out_0_19_1_port, P_OUT => 
                           lev_i_out_0_19_0_port);
   PG_NETWORK_0_20 : PG_NET_45 port map( A => A(19), B => B(19), G_OUT => 
                           lev_i_out_0_20_1_port, P_OUT => 
                           lev_i_out_0_20_0_port);
   PG_NETWORK_0_21 : PG_NET_44 port map( A => A(20), B => B(20), G_OUT => 
                           lev_i_out_0_21_1_port, P_OUT => 
                           lev_i_out_0_21_0_port);
   PG_NETWORK_0_22 : PG_NET_43 port map( A => A(21), B => B(21), G_OUT => 
                           lev_i_out_0_22_1_port, P_OUT => 
                           lev_i_out_0_22_0_port);
   PG_NETWORK_0_23 : PG_NET_42 port map( A => A(22), B => B(22), G_OUT => 
                           lev_i_out_0_23_1_port, P_OUT => 
                           lev_i_out_0_23_0_port);
   PG_NETWORK_0_24 : PG_NET_41 port map( A => A(23), B => B(23), G_OUT => 
                           lev_i_out_0_24_1_port, P_OUT => 
                           lev_i_out_0_24_0_port);
   PG_NETWORK_0_25 : PG_NET_40 port map( A => A(24), B => B(24), G_OUT => 
                           lev_i_out_0_25_1_port, P_OUT => 
                           lev_i_out_0_25_0_port);
   PG_NETWORK_0_26 : PG_NET_39 port map( A => A(25), B => B(25), G_OUT => 
                           lev_i_out_0_26_1_port, P_OUT => 
                           lev_i_out_0_26_0_port);
   PG_NETWORK_0_27 : PG_NET_38 port map( A => A(26), B => B(26), G_OUT => 
                           lev_i_out_0_27_1_port, P_OUT => 
                           lev_i_out_0_27_0_port);
   PG_NETWORK_0_28 : PG_NET_37 port map( A => A(27), B => B(27), G_OUT => 
                           lev_i_out_0_28_1_port, P_OUT => 
                           lev_i_out_0_28_0_port);
   PG_NETWORK_0_29 : PG_NET_36 port map( A => A(28), B => B(28), G_OUT => 
                           lev_i_out_0_29_1_port, P_OUT => 
                           lev_i_out_0_29_0_port);
   PG_NETWORK_0_30 : PG_NET_35 port map( A => A(29), B => B(29), G_OUT => 
                           lev_i_out_0_30_1_port, P_OUT => 
                           lev_i_out_0_30_0_port);
   PG_NETWORK_0_31 : PG_NET_34 port map( A => A(30), B => B(30), G_OUT => 
                           lev_i_out_0_31_1_port, P_OUT => 
                           lev_i_out_0_31_0_port);
   PG_NETWORK_0_32 : PG_NET_33 port map( A => A(31), B => B(31), G_OUT => 
                           lev_i_out_0_32_1_port, P_OUT => 
                           lev_i_out_0_32_0_port);
   PG_NETWORK_0_33 : PG_NET_32 port map( A => A(32), B => B(32), G_OUT => 
                           lev_i_out_0_33_1_port, P_OUT => 
                           lev_i_out_0_33_0_port, clk => clk);
   PG_NETWORK_0_34 : PG_NET_31 port map( A => A(33), B => B(33), G_OUT => 
                           lev_i_out_0_34_1_port, P_OUT => n30);
   PG_NETWORK_0_35 : PG_NET_30 port map( A => A(34), B => B(34), G_OUT => 
                           lev_i_out_0_35_1_port, P_OUT => 
                           lev_i_out_0_35_0_port);
   PG_NETWORK_0_36 : PG_NET_29 port map( A => A(35), B => B(35), G_OUT => 
                           lev_i_out_0_36_1_port, P_OUT => 
                           lev_i_out_0_36_0_port);
   PG_NETWORK_0_37 : PG_NET_28 port map( A => A(36), B => B(36), G_OUT => 
                           lev_i_out_0_37_1_port, P_OUT => 
                           lev_i_out_0_37_0_port);
   PG_NETWORK_0_38 : PG_NET_27 port map( A => A(37), B => B(37), G_OUT => 
                           lev_i_out_0_38_1_port, P_OUT => 
                           lev_i_out_0_38_0_port);
   PG_NETWORK_0_39 : PG_NET_26 port map( A => A(38), B => B(38), G_OUT => 
                           lev_i_out_0_39_1_port, P_OUT => 
                           lev_i_out_0_39_0_port);
   PG_NETWORK_0_40 : PG_NET_25 port map( A => A(39), B => B(39), G_OUT => 
                           lev_i_out_0_40_1_port, P_OUT => 
                           lev_i_out_0_40_0_port);
   PG_NETWORK_0_41 : PG_NET_24 port map( A => A(40), B => B(40), G_OUT => 
                           lev_i_out_0_41_1_port, P_OUT => 
                           lev_i_out_0_41_0_port);
   PG_NETWORK_0_42 : PG_NET_23 port map( A => A(41), B => B(41), G_OUT => 
                           lev_i_out_0_42_1_port, P_OUT => 
                           lev_i_out_0_42_0_port);
   PG_NETWORK_0_43 : PG_NET_22 port map( A => A(42), B => B(42), G_OUT => 
                           lev_i_out_0_43_1_port, P_OUT => 
                           lev_i_out_0_43_0_port);
   PG_NETWORK_0_44 : PG_NET_21 port map( A => A(43), B => B(43), G_OUT => 
                           lev_i_out_0_44_1_port, P_OUT => 
                           lev_i_out_0_44_0_port);
   PG_NETWORK_0_45 : PG_NET_20 port map( A => A(44), B => B(44), G_OUT => 
                           lev_i_out_0_45_1_port, P_OUT => 
                           lev_i_out_0_45_0_port);
   PG_NETWORK_0_46 : PG_NET_19 port map( A => A(45), B => B(45), G_OUT => 
                           lev_i_out_0_46_1_port, P_OUT => 
                           lev_i_out_0_46_0_port, clk => clk);
   GNET1_1_2 : G_GENERAL_0 port map( PG_ik(1) => net102722, PG_ik(0) => 
                           lev_i_out_0_2_0_port, G_k_1j => lev_i_out_0_1_1_port
                           , G_ij => n27);
   PGNET1_1_4 : PG_GENERAL_0 port map( PG_ik(1) => lev_i_out_0_4_1_port, 
                           PG_ik(0) => lev_i_out_0_4_0_port, PG_k_1j(1) => 
                           lev_i_out_0_3_1_port, PG_k_1j(0) => 
                           lev_i_out_0_3_0_port, PG_ij(1) => 
                           lev_i_out_1_4_1_port, PG_ij(0) => 
                           lev_i_out_1_4_0_port);
   PGNET1_1_6 : PG_GENERAL_79 port map( PG_ik(1) => lev_i_out_0_6_1_port, 
                           PG_ik(0) => lev_i_out_0_6_0_port, PG_k_1j(1) => 
                           lev_i_out_0_5_1_port, PG_k_1j(0) => 
                           lev_i_out_0_5_0_port, PG_ij(1) => 
                           lev_i_out_1_6_1_port, PG_ij(0) => 
                           lev_i_out_1_6_0_port);
   PGNET1_1_8 : PG_GENERAL_78 port map( PG_ik(1) => lev_i_out_0_8_1_port, 
                           PG_ik(0) => lev_i_out_0_8_0_port, PG_k_1j(1) => 
                           lev_i_out_0_7_1_port, PG_k_1j(0) => 
                           lev_i_out_0_7_0_port, PG_ij(1) => 
                           lev_i_out_1_8_1_port, PG_ij(0) => 
                           lev_i_out_1_8_0_port);
   PGNET1_1_10 : PG_GENERAL_77 port map( PG_ik(1) => lev_i_out_0_10_1_port, 
                           PG_ik(0) => lev_i_out_0_10_0_port, PG_k_1j(1) => 
                           lev_i_out_0_9_1_port, PG_k_1j(0) => 
                           lev_i_out_0_9_0_port, PG_ij(1) => 
                           lev_i_out_1_10_1_port, PG_ij(0) => 
                           lev_i_out_1_10_0_port);
   PGNET1_1_12 : PG_GENERAL_76 port map( PG_ik(1) => lev_i_out_0_12_1_port, 
                           PG_ik(0) => lev_i_out_0_12_0_port, PG_k_1j(1) => 
                           lev_i_out_0_11_1_port, PG_k_1j(0) => 
                           lev_i_out_0_11_0_port, PG_ij(1) => 
                           lev_i_out_1_12_1_port, PG_ij(0) => 
                           lev_i_out_1_12_0_port);
   PGNET1_1_14 : PG_GENERAL_75 port map( PG_ik(1) => lev_i_out_0_14_1_port, 
                           PG_ik(0) => lev_i_out_0_14_0_port, PG_k_1j(1) => 
                           lev_i_out_0_13_1_port, PG_k_1j(0) => 
                           lev_i_out_0_13_0_port, PG_ij(1) => 
                           lev_i_out_1_14_1_port, PG_ij(0) => 
                           lev_i_out_1_14_0_port);
   PGNET1_1_16 : PG_GENERAL_74 port map( PG_ik(1) => lev_i_out_0_16_1_port, 
                           PG_ik(0) => lev_i_out_0_16_0_port, PG_k_1j(1) => 
                           lev_i_out_0_15_1_port, PG_k_1j(0) => 
                           lev_i_out_0_15_0_port, PG_ij(1) => 
                           lev_i_out_1_16_1_port, PG_ij(0) => 
                           lev_i_out_1_16_0_port);
   PGNET1_1_18 : PG_GENERAL_73 port map( PG_ik(1) => lev_i_out_0_18_1_port, 
                           PG_ik(0) => lev_i_out_0_18_0_port, PG_k_1j(1) => 
                           lev_i_out_0_17_1_port, PG_k_1j(0) => 
                           lev_i_out_0_17_0_port, PG_ij(1) => 
                           lev_i_out_1_18_1_port, PG_ij(0) => 
                           lev_i_out_1_18_0_port);
   PGNET1_1_20 : PG_GENERAL_72 port map( PG_ik(1) => lev_i_out_0_20_1_port, 
                           PG_ik(0) => lev_i_out_0_20_0_port, PG_k_1j(1) => 
                           lev_i_out_0_19_1_port, PG_k_1j(0) => 
                           lev_i_out_0_19_0_port, PG_ij(1) => 
                           lev_i_out_1_20_1_port, PG_ij(0) => 
                           lev_i_out_1_20_0_port);
   PGNET1_1_22 : PG_GENERAL_71 port map( PG_ik(1) => lev_i_out_0_22_1_port, 
                           PG_ik(0) => lev_i_out_0_22_0_port, PG_k_1j(1) => 
                           lev_i_out_0_21_1_port, PG_k_1j(0) => 
                           lev_i_out_0_21_0_port, PG_ij(1) => 
                           lev_i_out_1_22_1_port, PG_ij(0) => 
                           lev_i_out_1_22_0_port);
   PGNET1_1_24 : PG_GENERAL_70 port map( PG_ik(1) => lev_i_out_0_24_1_port, 
                           PG_ik(0) => lev_i_out_0_24_0_port, PG_k_1j(1) => 
                           lev_i_out_0_23_1_port, PG_k_1j(0) => 
                           lev_i_out_0_23_0_port, PG_ij(1) => 
                           lev_i_out_1_24_1_port, PG_ij(0) => 
                           lev_i_out_1_24_0_port);
   PGNET1_1_26 : PG_GENERAL_69 port map( PG_ik(1) => lev_i_out_0_26_1_port, 
                           PG_ik(0) => lev_i_out_0_26_0_port, PG_k_1j(1) => 
                           lev_i_out_0_25_1_port, PG_k_1j(0) => 
                           lev_i_out_0_25_0_port, PG_ij(1) => 
                           lev_i_out_1_26_1_port, PG_ij(0) => 
                           lev_i_out_1_26_0_port);
   PGNET1_1_28 : PG_GENERAL_68 port map( PG_ik(1) => lev_i_out_0_28_1_port, 
                           PG_ik(0) => lev_i_out_0_28_0_port, PG_k_1j(1) => 
                           lev_i_out_0_27_1_port, PG_k_1j(0) => 
                           lev_i_out_0_27_0_port, PG_ij(1) => 
                           lev_i_out_1_28_1_port, PG_ij(0) => 
                           lev_i_out_1_28_0_port);
   PGNET1_1_30 : PG_GENERAL_67 port map( PG_ik(1) => lev_i_out_0_30_1_port, 
                           PG_ik(0) => lev_i_out_0_30_0_port, PG_k_1j(1) => 
                           lev_i_out_0_29_1_port, PG_k_1j(0) => 
                           lev_i_out_0_29_0_port, PG_ij(1) => 
                           lev_i_out_1_30_1_port, PG_ij(0) => 
                           lev_i_out_1_30_0_port, clk => clk);
   PGNET1_1_32 : PG_GENERAL_66 port map( PG_ik(1) => lev_i_out_0_32_1_port, 
                           PG_ik(0) => lev_i_out_0_32_0_port, PG_k_1j(1) => 
                           lev_i_out_0_31_1_port, PG_k_1j(0) => 
                           lev_i_out_0_31_0_port, PG_ij(1) => 
                           lev_i_out_1_32_1_port, PG_ij(0) => 
                           lev_i_out_1_32_0_port);
   PGNET1_1_34 : PG_GENERAL_65 port map( PG_ik(1) => lev_i_out_0_34_1_port, 
                           PG_ik(0) => n30, PG_k_1j(1) => lev_i_out_0_33_1_port
                           , PG_k_1j(0) => lev_i_out_0_33_0_port, PG_ij(1) => 
                           lev_i_out_1_34_1_port, PG_ij(0) => 
                           lev_i_out_1_34_0_port, clk => clk);
   PGNET1_1_36 : PG_GENERAL_64 port map( PG_ik(1) => lev_i_out_0_36_1_port, 
                           PG_ik(0) => lev_i_out_0_36_0_port, PG_k_1j(1) => 
                           lev_i_out_0_35_1_port, PG_k_1j(0) => 
                           lev_i_out_0_35_0_port, PG_ij(1) => 
                           lev_i_out_1_36_1_port, PG_ij(0) => 
                           lev_i_out_1_36_0_port, clk => clk);
   PGNET1_1_38 : PG_GENERAL_63 port map( PG_ik(1) => lev_i_out_0_38_1_port, 
                           PG_ik(0) => lev_i_out_0_38_0_port, PG_k_1j(1) => 
                           lev_i_out_0_37_1_port, PG_k_1j(0) => 
                           lev_i_out_0_37_0_port, PG_ij(1) => 
                           lev_i_out_1_38_1_port, PG_ij(0) => 
                           lev_i_out_1_38_0_port, clk => clk);
   PGNET1_1_40 : PG_GENERAL_62 port map( PG_ik(1) => lev_i_out_0_40_1_port, 
                           PG_ik(0) => lev_i_out_0_40_0_port, PG_k_1j(1) => 
                           lev_i_out_0_39_1_port, PG_k_1j(0) => 
                           lev_i_out_0_39_0_port, PG_ij(1) => 
                           lev_i_out_1_40_1_port, PG_ij(0) => 
                           lev_i_out_1_40_0_port, clk => clk);
   PGNET1_1_42 : PG_GENERAL_61 port map( PG_ik(1) => lev_i_out_0_42_1_port, 
                           PG_ik(0) => lev_i_out_0_42_0_port, PG_k_1j(1) => 
                           lev_i_out_0_41_1_port, PG_k_1j(0) => 
                           lev_i_out_0_41_0_port, PG_ij(1) => 
                           lev_i_out_1_42_1_port, PG_ij(0) => 
                           lev_i_out_1_42_0_port, clk => clk);
   PGNET1_1_44 : PG_GENERAL_60 port map( PG_ik(1) => lev_i_out_0_44_1_port, 
                           PG_ik(0) => lev_i_out_0_44_0_port, PG_k_1j(1) => 
                           lev_i_out_0_43_1_port, PG_k_1j(0) => 
                           lev_i_out_0_43_0_port, PG_ij(1) => 
                           lev_i_out_1_44_1_port, PG_ij(0) => 
                           lev_i_out_1_44_0_port, clk => clk);
   PGNET1_1_46 : PG_GENERAL_59 port map( PG_ik(1) => lev_i_out_0_46_1_port, 
                           PG_ik(0) => lev_i_out_0_46_0_port, PG_k_1j(1) => 
                           lev_i_out_0_45_1_port, PG_k_1j(0) => 
                           lev_i_out_0_45_0_port, PG_ij(1) => 
                           lev_i_out_1_46_1_port, PG_ij(0) => 
                           lev_i_out_1_46_0_port);
   GNET_i_2_4_0 : G_GENERAL_31 port map( PG_ik(1) => lev_i_out_1_4_1_port, 
                           PG_ik(0) => lev_i_out_1_4_0_port, G_k_1j => n27, 
                           G_ij => n26, clk => clk);
   PGNET_i_2_8_0 : PG_GENERAL_49 port map( PG_ik(1) => lev_i_out_1_8_1_port, 
                           PG_ik(0) => lev_i_out_1_8_0_port, PG_k_1j(1) => 
                           lev_i_out_1_6_1_port, PG_k_1j(0) => 
                           lev_i_out_1_6_0_port, PG_ij(1) => 
                           lev_i_out_2_8_1_port, PG_ij(0) => 
                           lev_i_out_2_8_0_port);
   PGNET_i_2_12_0 : PG_GENERAL_48 port map( PG_ik(1) => lev_i_out_1_12_1_port, 
                           PG_ik(0) => lev_i_out_1_12_0_port, PG_k_1j(1) => 
                           lev_i_out_1_10_1_port, PG_k_1j(0) => 
                           lev_i_out_1_10_0_port, PG_ij(1) => 
                           lev_i_out_2_12_1_port, PG_ij(0) => 
                           lev_i_out_2_12_0_port);
   PGNET_i_2_16_0 : PG_GENERAL_47 port map( PG_ik(1) => lev_i_out_1_16_1_port, 
                           PG_ik(0) => lev_i_out_1_16_0_port, PG_k_1j(1) => 
                           lev_i_out_1_14_1_port, PG_k_1j(0) => 
                           lev_i_out_1_14_0_port, PG_ij(1) => 
                           lev_i_out_2_16_1_port, PG_ij(0) => 
                           lev_i_out_2_16_0_port);
   PGNET_i_2_20_0 : PG_GENERAL_46 port map( PG_ik(1) => lev_i_out_1_20_1_port, 
                           PG_ik(0) => lev_i_out_1_20_0_port, PG_k_1j(1) => 
                           lev_i_out_1_18_1_port, PG_k_1j(0) => 
                           lev_i_out_1_18_0_port, PG_ij(1) => 
                           lev_i_out_2_20_1_port, PG_ij(0) => 
                           lev_i_out_2_20_0_port);
   PGNET_i_2_24_0 : PG_GENERAL_45 port map( PG_ik(1) => lev_i_out_1_24_1_port, 
                           PG_ik(0) => lev_i_out_1_24_0_port, PG_k_1j(1) => 
                           lev_i_out_1_22_1_port, PG_k_1j(0) => 
                           lev_i_out_1_22_0_port, PG_ij(1) => 
                           lev_i_out_2_24_1_port, PG_ij(0) => 
                           lev_i_out_2_24_0_port);
   PGNET_i_2_28_0 : PG_GENERAL_44 port map( PG_ik(1) => lev_i_out_1_28_1_port, 
                           PG_ik(0) => lev_i_out_1_28_0_port, PG_k_1j(1) => n23
                           , PG_k_1j(0) => n22, PG_ij(1) => 
                           lev_i_out_2_28_1_port, PG_ij(0) => 
                           lev_i_out_2_28_0_port, clk => clk);
   PGNET_i_2_32_0 : PG_GENERAL_43 port map( PG_ik(1) => lev_i_out_1_32_1_port, 
                           PG_ik(0) => lev_i_out_1_32_0_port, PG_k_1j(1) => 
                           lev_i_out_1_30_1_port, PG_k_1j(0) => n21, PG_ij(1) 
                           => lev_i_out_2_32_1_port, PG_ij(0) => 
                           lev_i_out_2_32_0_port, clk => clk);
   PGNET_i_2_36_0 : PG_GENERAL_42 port map( PG_ik(1) => lev_i_out_1_36_1_port, 
                           PG_ik(0) => lev_i_out_1_36_0_port, PG_k_1j(1) => 
                           lev_i_out_1_34_1_port, PG_k_1j(0) => 
                           lev_i_out_1_34_0_port, PG_ij(1) => 
                           lev_i_out_2_36_1_port, PG_ij(0) => 
                           lev_i_out_2_36_0_port);
   PGNET_i_2_40_0 : PG_GENERAL_41 port map( PG_ik(1) => lev_i_out_1_40_1_port, 
                           PG_ik(0) => lev_i_out_1_40_0_port, PG_k_1j(1) => 
                           lev_i_out_1_38_1_port, PG_k_1j(0) => 
                           lev_i_out_1_38_0_port, PG_ij(1) => 
                           lev_i_out_2_40_1_port, PG_ij(0) => 
                           lev_i_out_2_40_0_port);
   PGNET_i_2_44_0 : PG_GENERAL_40 port map( PG_ik(1) => lev_i_out_1_44_1_port, 
                           PG_ik(0) => lev_i_out_1_44_0_port, PG_k_1j(1) => 
                           lev_i_out_1_42_1_port, PG_k_1j(0) => 
                           lev_i_out_1_42_0_port, PG_ij(1) => 
                           lev_i_out_2_44_1_port, PG_ij(0) => 
                           lev_i_out_2_44_0_port);
   GNET_i_3_8_0 : G_GENERAL_29 port map( PG_ik(1) => lev_i_out_2_8_1_port, 
                           PG_ik(0) => lev_i_out_2_8_0_port, G_k_1j => n26, 
                           G_ij => n25);
   PGNET_i_3_16_0 : PG_GENERAL_33 port map( PG_ik(1) => lev_i_out_2_16_1_port, 
                           PG_ik(0) => lev_i_out_2_16_0_port, PG_k_1j(1) => 
                           lev_i_out_2_12_1_port, PG_k_1j(0) => 
                           lev_i_out_2_12_0_port, PG_ij(1) => 
                           lev_i_out_3_16_1_port, PG_ij(0) => 
                           lev_i_out_3_16_0_port);
   PGNET_i_3_22_2 : PG_GENERAL_32 port map( PG_ik(1) => lev_i_out_1_22_1_port, 
                           PG_ik(0) => lev_i_out_1_22_0_port, PG_k_1j(1) => n20
                           , PG_k_1j(0) => n19, PG_ij(1) => 
                           lev_i_out_3_22_1_port, PG_ij(0) => 
                           lev_i_out_3_22_0_port, clk => clk);
   PGNET_i_3_24_0 : PG_GENERAL_31 port map( PG_ik(1) => lev_i_out_2_24_1_port, 
                           PG_ik(0) => lev_i_out_2_24_0_port, PG_k_1j(1) => n20
                           , PG_k_1j(0) => n19, PG_ij(1) => n28, PG_ij(0) => 
                           lev_i_out_3_24_0_port, clk => clk);
   PGNET_i_3_30_2 : PG_GENERAL_30 port map( PG_ik(1) => lev_i_out_1_30_1_port, 
                           PG_ik(0) => n21, PG_k_1j(1) => lev_i_out_2_28_1_port
                           , PG_k_1j(0) => lev_i_out_2_28_0_port, PG_ij(1) => 
                           lev_i_out_3_30_1_port, PG_ij(0) => 
                           lev_i_out_3_30_0_port);
   PGNET_i_3_32_0 : PG_GENERAL_29 port map( PG_ik(1) => lev_i_out_2_32_1_port, 
                           PG_ik(0) => lev_i_out_2_32_0_port, PG_k_1j(1) => 
                           lev_i_out_2_28_1_port, PG_k_1j(0) => 
                           lev_i_out_2_28_0_port, PG_ij(1) => 
                           lev_i_out_3_32_1_port, PG_ij(0) => 
                           lev_i_out_3_32_0_port);
   PGNET_i_3_38_2 : PG_GENERAL_28 port map( PG_ik(1) => lev_i_out_1_38_1_port, 
                           PG_ik(0) => lev_i_out_1_38_0_port, PG_k_1j(1) => 
                           lev_i_out_2_36_1_port, PG_k_1j(0) => 
                           lev_i_out_2_36_0_port, PG_ij(1) => 
                           lev_i_out_3_38_1_port, PG_ij(0) => 
                           lev_i_out_3_38_0_port);
   PGNET_i_3_40_0 : PG_GENERAL_27 port map( PG_ik(1) => lev_i_out_2_40_1_port, 
                           PG_ik(0) => lev_i_out_2_40_0_port, PG_k_1j(1) => 
                           lev_i_out_2_36_1_port, PG_k_1j(0) => 
                           lev_i_out_2_36_0_port, PG_ij(1) => n38, PG_ij(0) => 
                           lev_i_out_3_40_0_port);
   PGNET_i_3_46_2 : PG_GENERAL_26 port map( PG_ik(1) => lev_i_out_1_46_1_port, 
                           PG_ik(0) => lev_i_out_1_46_0_port, PG_k_1j(1) => 
                           lev_i_out_2_44_1_port, PG_k_1j(0) => 
                           lev_i_out_2_44_0_port, PG_ij(1) => 
                           lev_i_out_3_46_1_port, PG_ij(0) => 
                           lev_i_out_3_46_0_port);
   GNET_i_4_16_0 : G_GENERAL_25 port map( PG_ik(1) => lev_i_out_3_16_1_port, 
                           PG_ik(0) => lev_i_out_3_16_0_port, G_k_1j => n25, 
                           G_ij => n17, clk => clk);
   PGNET_i_4_26_6 : PG_GENERAL_20 port map( PG_ik(1) => n23, PG_ik(0) => n22, 
                           PG_k_1j(1) => n28, PG_k_1j(0) => 
                           lev_i_out_3_24_0_port, PG_ij(1) => 
                           lev_i_out_4_26_1_port, PG_ij(0) => 
                           lev_i_out_4_26_0_port);
   PGNET_i_4_28_4 : PG_GENERAL_19 port map( PG_ik(1) => lev_i_out_2_28_1_port, 
                           PG_ik(0) => lev_i_out_2_28_0_port, PG_k_1j(1) => n28
                           , PG_k_1j(0) => lev_i_out_3_24_0_port, PG_ij(1) => 
                           lev_i_out_4_28_1_port, PG_ij(0) => 
                           lev_i_out_4_28_0_port);
   PGNET_i_4_30_2 : PG_GENERAL_18 port map( PG_ik(1) => lev_i_out_3_30_1_port, 
                           PG_ik(0) => lev_i_out_3_30_0_port, PG_k_1j(1) => n28
                           , PG_k_1j(0) => lev_i_out_3_24_0_port, PG_ij(1) => 
                           lev_i_out_4_30_1_port, PG_ij(0) => 
                           lev_i_out_4_30_0_port);
   PGNET_i_4_32_0 : PG_GENERAL_17 port map( PG_ik(1) => lev_i_out_3_32_1_port, 
                           PG_ik(0) => lev_i_out_3_32_0_port, PG_k_1j(1) => n28
                           , PG_k_1j(0) => lev_i_out_3_24_0_port, PG_ij(1) => 
                           lev_i_out_4_32_1_port, PG_ij(0) => 
                           lev_i_out_4_32_0_port);
   PGNET_i_4_42_6 : PG_GENERAL_16 port map( PG_ik(1) => lev_i_out_1_42_1_port, 
                           PG_ik(0) => lev_i_out_1_42_0_port, PG_k_1j(1) => n38
                           , PG_k_1j(0) => lev_i_out_3_40_0_port, PG_ij(1) => 
                           lev_i_out_4_42_1_port, PG_ij(0) => 
                           lev_i_out_4_42_0_port);
   PGNET_i_4_44_4 : PG_GENERAL_15 port map( PG_ik(1) => lev_i_out_2_44_1_port, 
                           PG_ik(0) => lev_i_out_2_44_0_port, PG_k_1j(1) => n38
                           , PG_k_1j(0) => lev_i_out_3_40_0_port, PG_ij(1) => 
                           lev_i_out_4_44_1_port, PG_ij(0) => 
                           lev_i_out_4_44_0_port);
   PGNET_i_4_46_2 : PG_GENERAL_14 port map( PG_ik(1) => lev_i_out_3_46_1_port, 
                           PG_ik(0) => lev_i_out_3_46_0_port, PG_k_1j(1) => n38
                           , PG_k_1j(0) => lev_i_out_3_40_0_port, PG_ij(1) => 
                           lev_i_out_4_46_1_port, PG_ij(0) => 
                           lev_i_out_4_46_0_port);
   GNET_i_5_22_10 : G_GENERAL_22 port map( PG_ik(1) => lev_i_out_3_22_1_port, 
                           PG_ik(0) => lev_i_out_3_22_0_port, G_k_1j => n17, 
                           G_ij => Co_11_port);
   GNET_i_5_24_8 : G_GENERAL_21 port map( PG_ik(1) => n28, PG_ik(0) => 
                           lev_i_out_3_24_0_port, G_k_1j => n17, G_ij => 
                           Co_12_port);
   GNET_i_5_26_6 : G_GENERAL_20 port map( PG_ik(1) => lev_i_out_4_26_1_port, 
                           PG_ik(0) => lev_i_out_4_26_0_port, G_k_1j => n17, 
                           G_ij => Co_13_port);
   GNET_i_5_28_4 : G_GENERAL_19 port map( PG_ik(1) => lev_i_out_4_28_1_port, 
                           PG_ik(0) => lev_i_out_4_28_0_port, G_k_1j => n17, 
                           G_ij => Co_14_port);
   GNET_i_5_30_2 : G_GENERAL_18 port map( PG_ik(1) => lev_i_out_4_30_1_port, 
                           PG_ik(0) => lev_i_out_4_30_0_port, G_k_1j => n17, 
                           G_ij => Co_15_port);
   GNET_i_5_32_0 : G_GENERAL_17 port map( PG_ik(1) => lev_i_out_4_32_1_port, 
                           PG_ik(0) => lev_i_out_4_32_0_port, G_k_1j => n17, 
                           G_ij => n16);
   GNET_i_6_34_30 : G_GENERAL_16 port map( PG_ik(1) => lev_i_out_1_34_1_port, 
                           PG_ik(0) => lev_i_out_1_34_0_port, G_k_1j => n16, 
                           G_ij => Co_17_port);
   GNET_i_6_36_28 : G_GENERAL_15 port map( PG_ik(1) => lev_i_out_2_36_1_port, 
                           PG_ik(0) => lev_i_out_2_36_0_port, G_k_1j => n16, 
                           G_ij => Co_18_port);
   GNET_i_6_38_26 : G_GENERAL_14 port map( PG_ik(1) => lev_i_out_3_38_1_port, 
                           PG_ik(0) => lev_i_out_3_38_0_port, G_k_1j => n16, 
                           G_ij => Co_19_port);
   GNET_i_6_40_24 : G_GENERAL_13 port map( PG_ik(1) => n38, PG_ik(0) => 
                           lev_i_out_3_40_0_port, G_k_1j => n16, G_ij => 
                           Co_20_port);
   GNET_i_6_42_22 : G_GENERAL_12 port map( PG_ik(1) => lev_i_out_4_42_1_port, 
                           PG_ik(0) => lev_i_out_4_42_0_port, G_k_1j => n16, 
                           G_ij => Co_21_port);
   GNET_i_6_44_20 : G_GENERAL_11 port map( PG_ik(1) => lev_i_out_4_44_1_port, 
                           PG_ik(0) => lev_i_out_4_44_0_port, G_k_1j => n16, 
                           G_ij => Co_22_port);
   GNET_i_6_46_18 : G_GENERAL_10 port map( PG_ik(1) => lev_i_out_4_46_1_port, 
                           PG_ik(0) => lev_i_out_4_46_0_port, G_k_1j => n16, 
                           G_ij => Co_23_port);
   MY_CLK_r_REG85_S2 : DFF_X1 port map( D => lev_i_out_1_30_0_port, CK => clk, 
                           Q => n21, QN => n_1471);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPround_SIG_width28_DW01_inc_1 is

   port( A : in std_logic_vector (24 downto 0);  SUM : out std_logic_vector (24
         downto 0));

end FPround_SIG_width28_DW01_inc_1;

architecture SYN_USE_DEFA_ARCH_NAME of FPround_SIG_width28_DW01_inc_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n6, n7, n11, n14, n15, n16, n17, n18, n19, n23, n26, n27, n28, 
      n29, n31, n35, n38, n40, n41, n50, n51, n52, n56, n57, n61, n62, n63, n68
      , n71, n72, n73, n74, n76, n80, n83, n84, n85, n86, n94, n95, n96, n97, 
      n101, n105, n106, n113, n115, n116, n122, n123, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n197, n198, 
      n199 : std_logic;

begin
   
   U154 : AND2_X1 port map( A1 => n28, A2 => n6, ZN => n181);
   U155 : XNOR2_X1 port map( A => n182, B => A(3), ZN => SUM(3));
   U156 : NAND2_X1 port map( A1 => n122, A2 => A(2), ZN => n182);
   U157 : XOR2_X1 port map( A => n183, B => A(5), Z => SUM(5));
   U158 : NOR2_X1 port map( A1 => n198, A2 => n113, ZN => n183);
   U159 : XOR2_X1 port map( A => n184, B => A(6), Z => SUM(6));
   U160 : NOR2_X1 port map( A1 => n198, A2 => n105, ZN => n184);
   U161 : XOR2_X1 port map( A => n185, B => A(7), Z => SUM(7));
   U162 : NOR2_X1 port map( A1 => n198, A2 => n101, ZN => n185);
   U163 : XNOR2_X1 port map( A => n186, B => A(9), ZN => SUM(9));
   U164 : NAND2_X1 port map( A1 => n94, A2 => A(8), ZN => n186);
   U165 : XNOR2_X1 port map( A => n187, B => A(11), ZN => SUM(11));
   U166 : NAND2_X1 port map( A1 => n94, A2 => n80, ZN => n187);
   U167 : XNOR2_X1 port map( A => n188, B => A(13), ZN => SUM(13));
   U168 : NAND2_X1 port map( A1 => n68, A2 => n94, ZN => n188);
   U169 : XNOR2_X1 port map( A => n189, B => A(14), ZN => SUM(14));
   U170 : NAND2_X1 port map( A1 => n61, A2 => n94, ZN => n189);
   U171 : XNOR2_X1 port map( A => n190, B => A(15), ZN => SUM(15));
   U172 : NAND2_X1 port map( A1 => n56, A2 => n94, ZN => n190);
   U173 : XNOR2_X1 port map( A => n191, B => A(17), ZN => SUM(17));
   U174 : NAND2_X1 port map( A1 => n199, A2 => A(16), ZN => n191);
   U175 : XNOR2_X1 port map( A => n192, B => A(19), ZN => SUM(19));
   U176 : NAND2_X1 port map( A1 => n1, A2 => n35, ZN => n192);
   U177 : XNOR2_X1 port map( A => n193, B => A(21), ZN => SUM(21));
   U178 : NAND2_X1 port map( A1 => n199, A2 => n23, ZN => n193);
   U179 : XNOR2_X1 port map( A => n194, B => A(23), ZN => SUM(23));
   U180 : NAND2_X1 port map( A1 => n11, A2 => n199, ZN => n194);
   U181 : INV_X1 port map( A => n95, ZN => n94);
   U183 : INV_X1 port map( A => n73, ZN => n74);
   U185 : NOR2_X1 port map( A1 => n19, A2 => n7, ZN => n6);
   U186 : NOR2_X1 port map( A1 => n41, A2 => n38, ZN => n35);
   U187 : NOR2_X1 port map( A1 => n86, A2 => n83, ZN => n80);
   U188 : NOR2_X1 port map( A1 => n29, A2 => n26, ZN => n23);
   U189 : INV_X1 port map( A => n28, ZN => n29);
   U190 : INV_X1 port map( A => n123, ZN => n122);
   U191 : NOR2_X1 port map( A1 => n74, A2 => n62, ZN => n61);
   U192 : NOR2_X1 port map( A1 => n74, A2 => n71, ZN => n68);
   U193 : NOR2_X1 port map( A1 => n17, A2 => n14, ZN => n11);
   U194 : NAND2_X1 port map( A1 => n28, A2 => n18, ZN => n17);
   U195 : INV_X1 port map( A => n19, ZN => n18);
   U197 : NAND2_X1 port map( A1 => n73, A2 => n51, ZN => n50);
   U198 : NOR2_X1 port map( A1 => n62, A2 => n52, ZN => n51);
   U199 : NAND2_X1 port map( A1 => A(14), A2 => A(15), ZN => n52);
   U200 : NOR2_X1 port map( A1 => n41, A2 => n31, ZN => n28);
   U201 : NAND2_X1 port map( A1 => A(18), A2 => A(19), ZN => n31);
   U203 : NAND2_X1 port map( A1 => A(10), A2 => A(11), ZN => n76);
   U204 : NOR2_X1 port map( A1 => n116, A2 => n123, ZN => n115);
   U205 : NAND2_X1 port map( A1 => A(2), A2 => A(3), ZN => n116);
   U206 : XOR2_X1 port map( A => n199, B => A(16), Z => SUM(16));
   U207 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n41);
   U208 : NAND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n86);
   U209 : XOR2_X1 port map( A => n84, B => n83, Z => SUM(10));
   U210 : NAND2_X1 port map( A1 => n94, A2 => n85, ZN => n84);
   U211 : INV_X1 port map( A => n86, ZN => n85);
   U212 : XOR2_X1 port map( A => n72, B => n71, Z => SUM(12));
   U213 : NAND2_X1 port map( A1 => n94, A2 => n73, ZN => n72);
   U216 : INV_X1 port map( A => n41, ZN => n40);
   U217 : XOR2_X1 port map( A => n27, B => n26, Z => SUM(20));
   U218 : NAND2_X1 port map( A1 => n1, A2 => n28, ZN => n27);
   U219 : XOR2_X1 port map( A => n15, B => n14, Z => SUM(22));
   U220 : NAND2_X1 port map( A1 => n199, A2 => n16, ZN => n15);
   U221 : INV_X1 port map( A => n17, ZN => n16);
   U222 : INV_X1 port map( A => A(18), ZN => n38);
   U223 : INV_X1 port map( A => A(20), ZN => n26);
   U224 : INV_X1 port map( A => A(10), ZN => n83);
   U225 : INV_X1 port map( A => A(22), ZN => n14);
   U226 : INV_X1 port map( A => A(12), ZN => n71);
   U227 : INV_X1 port map( A => A(4), ZN => n113);
   U228 : XOR2_X1 port map( A => n198, B => n113, Z => SUM(4));
   U229 : NAND2_X1 port map( A1 => A(4), A2 => A(5), ZN => n105);
   U230 : NAND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n62);
   U231 : XOR2_X1 port map( A => n94, B => A(8), Z => SUM(8));
   U232 : NOR2_X1 port map( A1 => n74, A2 => n57, ZN => n56);
   U233 : NAND2_X1 port map( A1 => n63, A2 => A(14), ZN => n57);
   U234 : INV_X1 port map( A => n62, ZN => n63);
   U235 : NAND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n123);
   U236 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n19);
   U237 : NAND2_X1 port map( A1 => n106, A2 => A(6), ZN => n101);
   U238 : INV_X1 port map( A => n105, ZN => n106);
   U239 : NAND2_X1 port map( A1 => A(22), A2 => A(23), ZN => n7);
   U240 : NAND2_X1 port map( A1 => n115, A2 => n96, ZN => n95);
   U241 : NOR2_X1 port map( A1 => n105, A2 => n97, ZN => n96);
   U242 : NAND2_X1 port map( A1 => A(6), A2 => A(7), ZN => n97);
   U243 : XOR2_X1 port map( A => n122, B => A(2), Z => SUM(2));
   U244 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U245 : XOR2_X1 port map( A => A(1), B => A(0), Z => SUM(1));
   U182 : NOR2_X1 port map( A1 => n86, A2 => n76, ZN => n73);
   U196 : AND2_X1 port map( A1 => n1, A2 => n181, ZN => SUM(24));
   U202 : XNOR2_X1 port map( A => n197, B => n38, ZN => SUM(18));
   U214 : AND2_X1 port map( A1 => n199, A2 => n40, ZN => n197);
   U215 : OR2_X1 port map( A1 => n116, A2 => n123, ZN => n198);
   U246 : NOR2_X1 port map( A1 => n50, A2 => n95, ZN => n199);
   U247 : NOR2_X1 port map( A1 => n50, A2 => n95, ZN => n1);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity P4_ADDER_NBIT64_NBIT_PER_BLOCK2_NBLOCKS32 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (63 downto 0);  Cout : out std_logic;  clk : in 
         std_logic);

end P4_ADDER_NBIT64_NBIT_PER_BLOCK2_NBLOCKS32;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT64_NBIT_PER_BLOCK2_NBLOCKS32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GENERATOR_NBIT_PER_BLOCK2_NBLOCKS32
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic_vector
            (31 downto 0);  S : out std_logic_vector (63 downto 0);  clk : in 
            std_logic);
   end component;
   
   component CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK2
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (32 downto 0);  clk : in std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n186, n187, carry_out_22_port, carry_out_21_port, carry_out_20_port, 
      carry_out_19_port, carry_out_18_port, carry_out_17_port, 
      carry_out_16_port, carry_out_15_port, carry_out_14_port, 
      carry_out_13_port, carry_out_12_port, carry_out_11_port, n5, n7, n14, n20
      , n21, n22, n29, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n171, n188, n189, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552,
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606 : 
      std_logic;

begin
   
   MY_CLK_r_REG219_S2 : DFF_X1 port map( D => A(44), CK => clk, Q => n14, QN =>
                           n_1546);
   MY_CLK_r_REG218_S2 : DFF_X1 port map( D => B(45), CK => clk, Q => n7, QN => 
                           n_1547);
   MY_CLK_r_REG209_S2 : DFF_X1 port map( D => B(44), CK => clk, Q => n5, QN => 
                           n_1548);
   n20 <= '0';
   n21 <= '0';
   n22 <= '0';
   n29 <= '0';
   n42 <= '0';
   n43 <= '0';
   n44 <= '0';
   n45 <= '0';
   n46 <= '0';
   n47 <= '0';
   n48 <= '0';
   n49 <= '0';
   n50 <= '0';
   n51 <= '0';
   n52 <= '0';
   n53 <= '0';
   n54 <= '0';
   n55 <= '0';
   n56 <= '0';
   n57 <= '0';
   n58 <= '0';
   n59 <= '0';
   n60 <= '0';
   n61 <= '0';
   n62 <= '0';
   n63 <= '0';
   n64 <= '0';
   n65 <= '0';
   n66 <= '0';
   n67 <= '0';
   n68 <= '0';
   n69 <= '0';
   n70 <= '0';
   n71 <= '0';
   n72 <= '0';
   n73 <= '0';
   n74 <= '0';
   n75 <= '0';
   n76 <= '0';
   n77 <= '0';
   n78 <= '0';
   n79 <= '0';
   n80 <= '0';
   n81 <= '0';
   n82 <= '0';
   n83 <= '0';
   n84 <= '0';
   n85 <= '0';
   n86 <= '0';
   n87 <= '0';
   n88 <= '0';
   n89 <= '0';
   n90 <= '0';
   n91 <= '0';
   n92 <= '0';
   n93 <= '0';
   n94 <= '0';
   n95 <= '0';
   n96 <= '0';
   n97 <= '0';
   n98 <= '0';
   n99 <= '0';
   n100 <= '0';
   n101 <= '0';
   n102 <= '0';
   n103 <= '0';
   n104 <= '0';
   n105 <= '0';
   n106 <= '0';
   n107 <= '0';
   n108 <= '0';
   n109 <= '0';
   n110 <= '0';
   n111 <= '0';
   n112 <= '0';
   n113 <= '0';
   n114 <= '0';
   n115 <= '0';
   n116 <= '0';
   n117 <= '0';
   n118 <= '0';
   n119 <= '0';
   n120 <= '0';
   n121 <= '0';
   n122 <= '0';
   n123 <= '0';
   n124 <= '0';
   n125 <= '0';
   n126 <= '0';
   n127 <= '0';
   n128 <= '0';
   n129 <= '0';
   n130 <= '0';
   n131 <= '0';
   n132 <= '0';
   n133 <= '0';
   n134 <= '0';
   n135 <= '0';
   n136 <= '0';
   n137 <= '0';
   n138 <= '0';
   n139 <= '0';
   n140 <= '0';
   n141 <= '0';
   n142 <= '0';
   n143 <= '0';
   n144 <= '0';
   n145 <= '0';
   n146 <= '0';
   n147 <= '0';
   n148 <= '0';
   n149 <= '0';
   n150 <= '0';
   n151 <= '0';
   n152 <= '0';
   n153 <= '0';
   n154 <= '0';
   n155 <= '0';
   n156 <= '0';
   n157 <= '0';
   n158 <= '0';
   n159 <= '0';
   n160 <= '0';
   n161 <= '0';
   n162 <= '0';
   n163 <= '0';
   n164 <= '0';
   n165 <= '0';
   n166 <= '0';
   n167 <= '0';
   n168 <= '0';
   n187 <= '0';
   n186 <= '0';
   CARRY_GEN_INST : CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK2 port map( A(63) => 
                           n20, A(62) => n21, A(61) => n22, A(60) => n29, A(59)
                           => n42, A(58) => n43, A(57) => n44, A(56) => n45, 
                           A(55) => n46, A(54) => n47, A(53) => n48, A(52) => 
                           n49, A(51) => n50, A(50) => n51, A(49) => n52, A(48)
                           => n53, A(47) => n54, A(46) => n55, A(45) => A(45), 
                           A(44) => n14, A(43) => A(43), A(42) => A(42), A(41) 
                           => A(41), A(40) => A(40), A(39) => A(39), A(38) => 
                           A(38), A(37) => A(37), A(36) => A(36), A(35) => 
                           A(35), A(34) => A(34), A(33) => A(33), A(32) => 
                           A(32), A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(63) => n56, B(62) => n57, B(61) => n58, 
                           B(60) => n59, B(59) => n60, B(58) => n61, B(57) => 
                           n62, B(56) => n63, B(55) => n64, B(54) => n65, B(53)
                           => n66, B(52) => n67, B(51) => n68, B(50) => n69, 
                           B(49) => n70, B(48) => n71, B(47) => n72, B(46) => 
                           n73, B(45) => n7, B(44) => n5, B(43) => B(43), B(42)
                           => B(42), B(41) => B(41), B(40) => B(40), B(39) => 
                           B(39), B(38) => B(38), B(37) => B(37), B(36) => 
                           B(36), B(35) => B(35), B(34) => B(34), B(33) => 
                           B(33), B(32) => B(32), B(31) => B(31), B(30) => 
                           B(30), B(29) => B(29), B(28) => B(28), B(27) => 
                           B(27), B(26) => B(26), B(25) => B(25), B(24) => 
                           B(24), B(23) => B(23), B(22) => B(22), B(21) => 
                           B(21), B(20) => B(20), B(19) => B(19), B(18) => 
                           B(18), B(17) => B(17), B(16) => B(16), B(15) => 
                           B(15), B(14) => B(14), B(13) => B(13), B(12) => 
                           B(12), B(11) => B(11), B(10) => B(10), B(9) => B(9),
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => n186, B(0) => B(0), Cin => n187, Co(32) => n_1549
                           , Co(31) => n_1550, Co(30) => n_1551, Co(29) => 
                           n_1552, Co(28) => n_1553, Co(27) => n_1554, Co(26) 
                           => n_1555, Co(25) => n_1556, Co(24) => n_1557, 
                           Co(23) => n171, Co(22) => carry_out_22_port, Co(21) 
                           => carry_out_21_port, Co(20) => carry_out_20_port, 
                           Co(19) => carry_out_19_port, Co(18) => 
                           carry_out_18_port, Co(17) => carry_out_17_port, 
                           Co(16) => carry_out_16_port, Co(15) => 
                           carry_out_15_port, Co(14) => carry_out_14_port, 
                           Co(13) => carry_out_13_port, Co(12) => 
                           carry_out_12_port, Co(11) => carry_out_11_port, 
                           Co(10) => n_1558, Co(9) => n_1559, Co(8) => n_1560, 
                           Co(7) => n_1561, Co(6) => n_1562, Co(5) => n_1563, 
                           Co(4) => n_1564, Co(3) => n_1565, Co(2) => n_1566, 
                           Co(1) => n_1567, Co(0) => n_1568, clk => clk);
   SUM_GEN_INST : SUM_GENERATOR_NBIT_PER_BLOCK2_NBLOCKS32 port map( A(63) => 
                           n74, A(62) => n75, A(61) => n76, A(60) => n77, A(59)
                           => n78, A(58) => n79, A(57) => n80, A(56) => n81, 
                           A(55) => n82, A(54) => n83, A(53) => n84, A(52) => 
                           n85, A(51) => n86, A(50) => n87, A(49) => n88, A(48)
                           => n89, A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => n14, A(43) => A(43), A(42) => A(42),
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => n188, A(32)
                           => A(32), A(31) => n189, A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => n90, A(20) => n91, 
                           A(19) => n92, A(18) => n93, A(17) => n94, A(16) => 
                           n95, A(15) => n96, A(14) => n97, A(13) => n98, A(12)
                           => n99, A(11) => n100, A(10) => n101, A(9) => n102, 
                           A(8) => n103, A(7) => n104, A(6) => n105, A(5) => 
                           n106, A(4) => n107, A(3) => n108, A(2) => n109, A(1)
                           => n110, A(0) => n111, B(63) => n112, B(62) => n113,
                           B(61) => n114, B(60) => n115, B(59) => n116, B(58) 
                           => n117, B(57) => n118, B(56) => n119, B(55) => n120
                           , B(54) => n121, B(53) => n122, B(52) => n123, B(51)
                           => n124, B(50) => n125, B(49) => n126, B(48) => n127
                           , B(47) => B(47), B(46) => B(46), B(45) => n7, B(44)
                           => n5, B(43) => B(43), B(42) => B(42), B(41) => 
                           B(41), B(40) => B(40), B(39) => B(39), B(38) => 
                           B(38), B(37) => B(37), B(36) => B(36), B(35) => 
                           B(35), B(34) => B(34), B(33) => B(33), B(32) => 
                           B(32), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => n128, B(20) => n129,
                           B(19) => n130, B(18) => n131, B(17) => n132, B(16) 
                           => n133, B(15) => n134, B(14) => n135, B(13) => n136
                           , B(12) => n137, B(11) => n138, B(10) => n139, B(9) 
                           => n140, B(8) => n141, B(7) => n142, B(6) => n143, 
                           B(5) => n144, B(4) => n145, B(3) => n146, B(2) => 
                           n147, B(1) => n148, B(0) => n149, Ci(31) => n150, 
                           Ci(30) => n151, Ci(29) => n152, Ci(28) => n153, 
                           Ci(27) => n154, Ci(26) => n155, Ci(25) => n156, 
                           Ci(24) => n157, Ci(23) => n171, Ci(22) => 
                           carry_out_22_port, Ci(21) => carry_out_21_port, 
                           Ci(20) => carry_out_20_port, Ci(19) => 
                           carry_out_19_port, Ci(18) => carry_out_18_port, 
                           Ci(17) => carry_out_17_port, Ci(16) => 
                           carry_out_16_port, Ci(15) => carry_out_15_port, 
                           Ci(14) => carry_out_14_port, Ci(13) => 
                           carry_out_13_port, Ci(12) => carry_out_12_port, 
                           Ci(11) => carry_out_11_port, Ci(10) => n158, Ci(9) 
                           => n159, Ci(8) => n160, Ci(7) => n161, Ci(6) => n162
                           , Ci(5) => n163, Ci(4) => n164, Ci(3) => n165, Ci(2)
                           => n166, Ci(1) => n167, Ci(0) => n168, S(63) => 
                           n_1569, S(62) => n_1570, S(61) => n_1571, S(60) => 
                           n_1572, S(59) => n_1573, S(58) => n_1574, S(57) => 
                           n_1575, S(56) => n_1576, S(55) => n_1577, S(54) => 
                           n_1578, S(53) => n_1579, S(52) => n_1580, S(51) => 
                           n_1581, S(50) => n_1582, S(49) => n_1583, S(48) => 
                           n_1584, S(47) => S(47), S(46) => S(46), S(45) => 
                           S(45), S(44) => S(44), S(43) => S(43), S(42) => 
                           S(42), S(41) => S(41), S(40) => S(40), S(39) => 
                           S(39), S(38) => S(38), S(37) => S(37), S(36) => 
                           S(36), S(35) => S(35), S(34) => S(34), S(33) => 
                           S(33), S(32) => S(32), S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           n_1585, S(20) => n_1586, S(19) => n_1587, S(18) => 
                           n_1588, S(17) => n_1589, S(16) => n_1590, S(15) => 
                           n_1591, S(14) => n_1592, S(13) => n_1593, S(12) => 
                           n_1594, S(11) => n_1595, S(10) => n_1596, S(9) => 
                           n_1597, S(8) => n_1598, S(7) => n_1599, S(6) => 
                           n_1600, S(5) => n_1601, S(4) => n_1602, S(3) => 
                           n_1603, S(2) => n_1604, S(1) => n_1605, S(0) => 
                           n_1606, clk => clk);
   U4 : CLKBUF_X1 port map( A => A(33), Z => n188);
   U6 : BUF_X1 port map( A => A(31), Z => n189);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U2 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U1 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U2 : XOR2_X1 port map( A => A, B => B, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_153 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n3, B => n1, ZN => S);
   U1 : INV_X1 port map( A => A, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n1, A2 => B_BAR, ZN => Co);
   U4 : INV_X1 port map( A => B_BAR, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U4 : XOR2_X1 port map( A => A, B => B, Z => S);
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U1 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => Co);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n3);
   U1 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => Co);
   U2 : XOR2_X1 port map( A => A, B => B, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29785, net29786, net29787, n1, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => n4, B2 => B, A => Ci, ZN => net29787);
   U4 : INV_X1 port map( A => B, ZN => net29786);
   U6 : INV_X1 port map( A => n4, ZN => net29785);
   U7 : OAI21_X1 port map( B1 => net29785, B2 => net29786, A => net29787, ZN =>
                           Co);
   U5 : CLKBUF_X1 port map( A => A, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n7);
   U7 : XNOR2_X1 port map( A => A, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   U2 : XNOR2_X1 port map( A => n5, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n7 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U5 : INV_X1 port map( A => n7, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n3);
   U7 : OAI21_X1 port map( B1 => n7, B2 => B, A => Ci, ZN => n2);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : CLKBUF_X1 port map( A => A, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => n7, ZN => S);
   U2 : NAND2_X1 port map( A1 => n8, A2 => Ci, ZN => n3);
   U3 : NAND2_X1 port map( A1 => A, A2 => n1, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : INV_X1 port map( A => A, ZN => n8);
   U8 : INV_X1 port map( A => B, ZN => n7);
   U9 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n6);
   U10 : OAI21_X1 port map( B1 => n8, B2 => n7, A => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U1 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n3);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => B, Z => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG405_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG418_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n_1617 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n6, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => n6, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG464_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1617);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5, n7, n9 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n7, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n9, B1 => n3, B2 => n2, ZN => Co);
   MY_CLK_r_REG423_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n9)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG462_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   MY_CLK_r_REG455_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG461_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n11, B1 => n2, B2 => n10, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => n8, ZN => n4);
   MY_CLK_r_REG493_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );
   MY_CLK_r_REG402_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n13, n_1618 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n10, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG403_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1618);
   MY_CLK_r_REG473_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   MY_CLK_r_REG421_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n13, n_1619 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n10, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG422_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1619);
   MY_CLK_r_REG494_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   MY_CLK_r_REG438_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_204 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => Ci_BAR, A2 => n4, B1 => n2, B2 => n1, ZN => Co
                           );
   U3 : INV_X1 port map( A => Ci_BAR, ZN => n6);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_205 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => n2, B2 => n1, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_206 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n1, A2 => n6, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29953, net29954, net29955, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net29955);
   U4 : INV_X1 port map( A => A, ZN => net29953);
   U5 : INV_X1 port map( A => B, ZN => net29954);
   U7 : OAI21_X1 port map( B1 => net29953, B2 => net29954, A => net29955, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co_BAR : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n1);
   U4 : AND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U5 : OAI22_X1 port map( A1 => n2, A2 => n3, B1 => Ci, B2 => n3, ZN => Co_BAR
                           );
   U3 : XNOR2_X1 port map( A => A, B => n6, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29979, net29980, net29981, n1, n3 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n1);
   U3 : XNOR2_X1 port map( A => n1, B => Ci, ZN => S);
   U4 : INV_X1 port map( A => B, ZN => net29980);
   U5 : OAI21_X1 port map( B1 => n3, B2 => B, A => Ci, ZN => net29981);
   U7 : INV_X1 port map( A => n3, ZN => net29979);
   U8 : OAI21_X1 port map( B1 => net29979, B2 => net29980, A => net29981, ZN =>
                           Co);
   U1 : CLKBUF_X1 port map( A => A, Z => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => A, ZN => n3);
   U7 : INV_X1 port map( A => B, ZN => n2);
   U1 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U5 : INV_X1 port map( A => n1, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => n8, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n6);
   U4 : XNOR2_X1 port map( A => n6, B => A, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U8 : INV_X1 port map( A => Ci, ZN => n2);
   U1 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n7 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => n7, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n6);
   U4 : XNOR2_X1 port map( A => A, B => n6, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U8 : INV_X1 port map( A => Ci, ZN => n2);
   U2 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n7 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n7);
   U2 : XNOR2_X1 port map( A => A, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U1 : XNOR2_X1 port map( A => n7, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n1);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U4 : OAI22_X1 port map( A1 => n2, A2 => n1, B1 => Ci, B2 => n2, ZN => n4);
   U5 : INV_X1 port map( A => n4, ZN => Co);
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => n2, ZN => n5);
   U3 : AND2_X1 port map( A1 => Ci, A2 => n6, ZN => n2);
   U4 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U6 : INV_X1 port map( A => A, ZN => n7);
   U7 : INV_X1 port map( A => B, ZN => n6);
   U8 : INV_X1 port map( A => Ci, ZN => n3);
   U9 : NOR2_X1 port map( A1 => n3, A2 => A, ZN => n4);
   U10 : OAI21_X1 port map( B1 => n7, B2 => n6, A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => n2, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U5 : XNOR2_X1 port map( A => n6, B => n5, ZN => n8);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U7 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n6);
   U8 : INV_X1 port map( A => A, ZN => n3);
   U9 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => Co);
   U10 : INV_X1 port map( A => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => n6, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n6, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n8, A => n1, ZN => Co);
   MY_CLK_r_REG329_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => n6, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n6, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n8, A => n1, ZN => Co);
   MY_CLK_r_REG342_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n10, B2 => n11, ZN => Co);
   MY_CLK_r_REG349_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n11)
                           ;
   MY_CLK_r_REG343_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n10)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n14, B1 => n12, B2 => n13, ZN => Co)
                           ;
   MY_CLK_r_REG406_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n14
                           );
   MY_CLK_r_REG359_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG350_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6, n7, n_1621, n_1622 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => n6, B => n7, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => n7, A => n6, ZN => n3);
   MY_CLK_r_REG371_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => 
                           n_1621);
   MY_CLK_r_REG419_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1622);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1623, n_1624 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG372_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1623, QN => 
                           n13);
   MY_CLK_r_REG378_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1624, QN => 
                           n14);
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);
   MY_CLK_r_REG465_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n14, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG424_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   MY_CLK_r_REG383_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG379_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n14
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n14, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG463_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   MY_CLK_r_REG389_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG384_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n14
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n9, n10, n11, n12, n14, n_1625, n_1626, n_1627 : 
      std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n9, A2 => n14, B1 => n12, B2 => n11, ZN => Co)
                           ;
   MY_CLK_r_REG390_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n12, QN => 
                           n_1625);
   MY_CLK_r_REG394_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n11, QN => 
                           n_1626);
   MY_CLK_r_REG391_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n9, QN => 
                           n_1627);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   MY_CLK_r_REG454_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1628 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG404_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1628, QN => 
                           n14);
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);
   MY_CLK_r_REG460_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   MY_CLK_r_REG395_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n8, n_1630, n_1631 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => n8, B => n5, Z => n4);
   MY_CLK_r_REG231_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1630, QN => 
                           n8);
   MY_CLK_r_REG296_S1 : DFF_X1 port map( D => B, CK => clk, Q => n5, QN => 
                           n_1631);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  Co, S_BAR : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => S_BAR);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_258 is

   port( A, Ci : in std_logic;  Co : out std_logic;  B_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n6 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => n6, Z => S_BAR);
   U1 : INV_X1 port map( A => B_BAR, ZN => n6);
   U4 : NOR2_X1 port map( A1 => n2, A2 => B_BAR, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_259 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U1 : XNOR2_X1 port map( A => n2, B => n7, ZN => S);
   U3 : INV_X1 port map( A => B_BAR, ZN => n7);
   U4 : NOR2_X1 port map( A1 => n2, A2 => B_BAR, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_260 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U1 : NOR2_X1 port map( A1 => n2, A2 => B_BAR, ZN => Co);
   U3 : XNOR2_X1 port map( A => n2, B => n7, ZN => S);
   U4 : INV_X1 port map( A => B_BAR, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  Co, S : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n_1642 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n6, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => n6, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG415_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1642);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1643 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG411_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1643);
   MY_CLK_r_REG414_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => n6, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n8, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG324_S1 : DFF_X1 port map( D => A, CK => clk, Q => n6, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => n6, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => n6, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n8, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG293_S1 : DFF_X1 port map( D => A, CK => clk, Q => n6, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n7, n8, n10, n_1644 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => n8, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG409_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1644);
   MY_CLK_r_REG322_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n10)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => n8, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n11, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n10, B => n11, ZN => n4);
   MY_CLK_r_REG431_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n10
                           );
   MY_CLK_r_REG318_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n11)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n13, n_1645 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n10, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG320_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1645);
   MY_CLK_r_REG433_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   MY_CLK_r_REG432_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n8, n9, n12, n13 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U6 : OAI21_X1 port map( B1 => n9, B2 => A, A => n8, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n13, A => n2, ZN => Co);
   MY_CLK_r_REG434_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG440_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XNOR2_X1 port map( A => n12, B => n13, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n5, n9, n10, n11, n13, n14, n_1646 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n10, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => n9, B => n11, ZN => n5);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n11, A => n9, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n14, B2 => n13, A => n2, ZN => Co);
   MY_CLK_r_REG352_S1 : DFF_X1 port map( D => A, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG441_S1 : DFF_X1 port map( D => B, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG429_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => 
                           n_1646);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1647, n_1648 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG360_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1647, QN => 
                           n13);
   MY_CLK_r_REG430_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1648, QN => 
                           n14);
   MY_CLK_r_REG471_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1649, n_1650 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG373_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1649, QN => 
                           n13);
   MY_CLK_r_REG472_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1650, QN => 
                           n14);
   MY_CLK_r_REG427_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1651 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG399_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG428_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1651, QN => 
                           n14);
   MY_CLK_r_REG469_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n13, n_1652 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n13, ZN => Co)
                           ;
   MY_CLK_r_REG380_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1652);
   MY_CLK_r_REG470_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG425_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1653 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG398_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG426_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1653, QN => 
                           n14);
   MY_CLK_r_REG467_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1654 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG392_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG468_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1654, QN => 
                           n14);
   MY_CLK_r_REG457_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n9, n10, n11, n12, n14, n_1655, n_1656, n_1657 : 
      std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n9, A2 => n14, B1 => n12, B2 => n11, ZN => Co)
                           ;
   MY_CLK_r_REG396_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n12, QN => 
                           n_1655);
   MY_CLK_r_REG456_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n11, QN => 
                           n_1656);
   MY_CLK_r_REG466_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n14);
   MY_CLK_r_REG397_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n9, QN => 
                           n_1657);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_290 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => n2, B2 => n1, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n5, n6, n_1659, n_1660 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => n4, ZN => S);
   MY_CLK_r_REG229_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => 
                           n_1659);
   MY_CLK_r_REG228_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n5, QN => 
                           n_1660);
   U2 : XNOR2_X1 port map( A => A, B => n6, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n7, n10, n11, n_1661 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => n10, B => n7, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n10, B2 => n11, ZN => Co);
   MY_CLK_r_REG230_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1661, QN => 
                           n10);
   MY_CLK_r_REG233_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n11)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n8, n_1662 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : XOR2_X1 port map( A => n8, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n8, B2 => n1, ZN => Co);
   MY_CLK_r_REG234_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1662, QN => 
                           n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => n6, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n8, ZN => Co);
   MY_CLK_r_REG479_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U5 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net30323, net30324, net30325, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => net30323);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net30325);
   U5 : INV_X1 port map( A => B, ZN => net30324);
   U6 : OAI21_X1 port map( B1 => net30323, B2 => net30324, A => net30325, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => A, ZN => n2);
   U7 : INV_X1 port map( A => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_317;

architecture SYN_BEHAVIORAL of FA_317 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_318;

architecture SYN_BEHAVIORAL of FA_318 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : INV_X1 port map( A => Ci, ZN => n2);
   U3 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_319;

architecture SYN_BEHAVIORAL of FA_319 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net30350, net30351, net30352, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => B, ZN => net30351);
   U4 : INV_X1 port map( A => A, ZN => net30350);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net30352);
   U8 : OAI21_X1 port map( B1 => net30350, B2 => net30351, A => net30352, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_320;

architecture SYN_BEHAVIORAL of FA_320 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_321;

architecture SYN_BEHAVIORAL of FA_321 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n9 : std_logic;

begin
   
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => A, ZN => n4);
   U8 : INV_X1 port map( A => B, ZN => n3);
   U9 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);
   U1 : XNOR2_X1 port map( A => n9, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_322;

architecture SYN_BEHAVIORAL of FA_322 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n8, n9 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => B, B => n6, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => A, ZN => n6);
   U1 : NAND2_X2 port map( A1 => n9, A2 => n8, ZN => Co);
   U2 : NAND2_X2 port map( A1 => A, A2 => B, ZN => n8);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_323;

architecture SYN_BEHAVIORAL of FA_323 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_324;

architecture SYN_BEHAVIORAL of FA_324 is

   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => n7);
   U8 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n8);
   U9 : AND2_X2 port map( A1 => n7, A2 => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_325;

architecture SYN_BEHAVIORAL of FA_325 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => Co);
   U2 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U5 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U6 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_326;

architecture SYN_BEHAVIORAL of FA_326 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => A, ZN => n4);
   U8 : INV_X1 port map( A => B, ZN => n3);
   U9 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_327;

architecture SYN_BEHAVIORAL of FA_327 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7, n10, n11, n13, n14 : std_logic;

begin
   
   U4 : XNOR2_X1 port map( A => n7, B => n10, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => n11, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n11, A2 => A, ZN => n6);
   U8 : INV_X1 port map( A => A, ZN => n4);
   MY_CLK_r_REG100_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n13
                           );
   MY_CLK_r_REG323_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n14);
   U2 : AOI22_X1 port map( A1 => n6, A2 => n14, B1 => n4, B2 => n13, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_328;

architecture SYN_BEHAVIORAL of FA_328 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1663 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U2 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n1, ZN => Co);
   MY_CLK_r_REG101_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG110_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG319_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1663);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_329;

architecture SYN_BEHAVIORAL of FA_329 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n14, A => n1, ZN => Co);
   MY_CLK_r_REG111_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG267_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG321_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_330;

architecture SYN_BEHAVIORAL of FA_330 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n10, n11, n12, n14, n15, n16 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n11, B => n6, ZN => S);
   U3 : XNOR2_X1 port map( A => n12, B => n10, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => n5);
   U8 : AOI22_X1 port map( A1 => n5, A2 => n16, B1 => n15, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG265_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n15
                           );
   MY_CLK_r_REG275_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG339_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n16);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_331;

architecture SYN_BEHAVIORAL of FA_331 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n5, n9, n10, n11, n13, n14, n15 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n10, B => n5, ZN => S);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n11, A => n9, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n15, B2 => n13, A => n2, ZN => Co);
   MY_CLK_r_REG276_S1 : DFF_X1 port map( D => A, CK => clk, Q => n11, QN => n15
                           );
   MY_CLK_r_REG290_S1 : DFF_X1 port map( D => B, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG353_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => n14
                           );
   U1 : XNOR2_X1 port map( A => n14, B => n15, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_332;

architecture SYN_BEHAVIORAL of FA_332 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5, n8, n9, n11, n_1664 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n2, B => n9, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => n8, ZN => n2);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U6 : OAI21_X1 port map( B1 => n9, B2 => A, A => n8, ZN => n3);
   U7 : OAI21_X1 port map( B1 => n5, B2 => n11, A => n3, ZN => Co);
   MY_CLK_r_REG298_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n11)
                           ;
   MY_CLK_r_REG361_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1664);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_333;

architecture SYN_BEHAVIORAL of FA_333 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n7, n8, n10, n_1665 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U5 : OAI21_X1 port map( B1 => A, B2 => n8, A => n7, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n10, A => n2, ZN => Co);
   MY_CLK_r_REG306_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG374_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1665);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_334;

architecture SYN_BEHAVIORAL of FA_334 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n_1666, n_1667, n_1668 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n8, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => n7, B => n9, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n3);
   MY_CLK_r_REG307_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1666);
   MY_CLK_r_REG316_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1667);
   MY_CLK_r_REG400_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1668);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_335;

architecture SYN_BEHAVIORAL of FA_335 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1669 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n8, B => n9, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n13, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG317_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG327_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG381_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1669);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_336;

architecture SYN_BEHAVIORAL of FA_336 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6, n7, n_1670, n_1671 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   MY_CLK_r_REG328_S1 : DFF_X1 port map( D => A, CK => clk, Q => n7, QN => 
                           n_1670);
   MY_CLK_r_REG341_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n6, QN => 
                           n_1671);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_338;

architecture SYN_BEHAVIORAL of FA_338 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_339;

architecture SYN_BEHAVIORAL of FA_339 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n9, n_1672, n_1673 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => Ci, B => B, Z => n3);
   MY_CLK_r_REG358_S1 : DFF_X1 port map( D => A, CK => clk, Q => n7, QN => 
                           n_1672);
   MY_CLK_r_REG370_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n_1673, QN =>
                           n9);
   U5 : XNOR2_X1 port map( A => n7, B => n9, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_341;

architecture SYN_BEHAVIORAL of FA_341 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_342;

architecture SYN_BEHAVIORAL of FA_342 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_11 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_11;

architecture SYN_rtl of HA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_349 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_349;

architecture SYN_BEHAVIORAL of FA_349 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_350 is

   port( A : in std_logic;  S, Co : out std_logic;  clk, Ci_BAR, B_BAR : in 
         std_logic);

end FA_350;

architecture SYN_BEHAVIORAL of FA_350 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n7, n9, n_1675 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U5 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n7, B2 => B_BAR, ZN =>
                           Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => n9, B => n5, Z => S);
   MY_CLK_r_REG310_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n7, QN => 
                           n_1675);
   U2 : INV_X1 port map( A => Ci_BAR, ZN => n9);
   U3 : XNOR2_X1 port map( A => n7, B => B_BAR, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_363 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_363;

architecture SYN_BEHAVIORAL of FA_363 is

begin
   S <= B;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_364 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  clk, A_BAR : in 
         std_logic);

end FA_364;

architecture SYN_BEHAVIORAL of FA_364 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n6, n_1680 : std_logic;

begin
   
   U4 : INV_X1 port map( A => n6, ZN => n2);
   MY_CLK_r_REG416_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => 
                           n_1680);
   U1 : NOR2_X1 port map( A1 => A_BAR, A2 => n2, ZN => Co);
   U2 : XNOR2_X1 port map( A => A_BAR, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_365 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  clk, B_BAR : in 
         std_logic);

end FA_365;

architecture SYN_BEHAVIORAL of FA_365 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => B_BAR, ZN => S);
   MY_CLK_r_REG417_S1 : DFF_X1 port map( D => A, CK => clk, Q => n6, QN => n8);
   U2 : NOR2_X1 port map( A1 => n8, A2 => B_BAR, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_366;

architecture SYN_BEHAVIORAL of FA_366 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n_1683 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => n1, ZN => S);
   MY_CLK_r_REG413_S1 : DFF_X1 port map( D => B, CK => clk, Q => n5, QN => 
                           n_1683);
   U2 : AND2_X1 port map( A1 => A, A2 => n5, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_367;

architecture SYN_BEHAVIORAL of FA_367 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_368;

architecture SYN_BEHAVIORAL of FA_368 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n7, n8, n_1685, n_1686 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   MY_CLK_r_REG410_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1685);
   MY_CLK_r_REG445_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1686);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_369;

architecture SYN_BEHAVIORAL of FA_369 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1687 : std_logic;

begin
   
   U3 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n13, B2 => n12, A => n1, ZN => Co);
   U5 : XOR2_X1 port map( A => n8, B => n9, Z => n4);
   MY_CLK_r_REG412_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG443_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG475_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1687);
   U1 : XNOR2_X1 port map( A => n13, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_370;

architecture SYN_BEHAVIORAL of FA_370 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n8, n10, n11 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n8, B => n1, Z => S);
   MY_CLK_r_REG444_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n11)
                           ;
   MY_CLK_r_REG407_S1 : DFF_X1 port map( D => B, CK => clk, Q => n1, QN => n10)
                           ;
   U2 : NOR2_X1 port map( A1 => n11, A2 => n10, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_371;

architecture SYN_BEHAVIORAL of FA_371 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n_1689, n_1690 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => B, B => Ci, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   MY_CLK_r_REG408_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1689, QN => 
                           n9);
   MY_CLK_r_REG442_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n_1690, QN =>
                           n10);
   U1 : XOR2_X1 port map( A => n9, B => n10, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_372;

architecture SYN_BEHAVIORAL of FA_372 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_374;

architecture SYN_BEHAVIORAL of FA_374 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_387;

architecture SYN_BEHAVIORAL of FA_387 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_388 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_388;

architecture SYN_BEHAVIORAL of FA_388 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1693, n_1694 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG285_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1693);
   MY_CLK_r_REG232_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1694);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_389 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_389;

architecture SYN_BEHAVIORAL of FA_389 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1695 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG223_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG286_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1695, QN => 
                           n14);
   MY_CLK_r_REG273_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_390 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_390;

architecture SYN_BEHAVIORAL of FA_390 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1696, n_1697 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG478_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1696, QN => 
                           n13);
   MY_CLK_r_REG274_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1697, QN => 
                           n14);
   MY_CLK_r_REG226_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_391;

architecture SYN_BEHAVIORAL of FA_391 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n13, n_1698 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n10, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG214_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1698);
   MY_CLK_r_REG227_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG271_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_392;

architecture SYN_BEHAVIORAL of FA_392 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1699 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG221_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG272_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1699, QN => 
                           n14);
   MY_CLK_r_REG283_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_393;

architecture SYN_BEHAVIORAL of FA_393 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n11, n12, n_1700 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n1, ZN => S);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n3);
   MY_CLK_r_REG208_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG284_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1700);
   MY_CLK_r_REG291_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );
   U2 : XNOR2_X1 port map( A => n11, B => n12, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_394;

architecture SYN_BEHAVIORAL of FA_394 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1701 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG194_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG292_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1701, QN => 
                           n14);
   MY_CLK_r_REG303_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_395;

architecture SYN_BEHAVIORAL of FA_395 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1702 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n8, B => n10, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n1, ZN => Co);
   MY_CLK_r_REG204_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG304_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG308_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1702);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_396;

architecture SYN_BEHAVIORAL of FA_396 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n14, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG179_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n14
                           );
   MY_CLK_r_REG309_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG332_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_397;

architecture SYN_BEHAVIORAL of FA_397 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n10, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n1, ZN => Co);
   MY_CLK_r_REG192_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG333_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG311_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n14
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_398;

architecture SYN_BEHAVIORAL of FA_398 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n5, n9, n10, n11, n13, n14, n15 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => n11, ZN => S);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n11, A => n9, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n13, B2 => n14, A => n2, ZN => Co);
   MY_CLK_r_REG164_S1 : DFF_X1 port map( D => A, CK => clk, Q => n11, QN => n13
                           );
   MY_CLK_r_REG312_S1 : DFF_X1 port map( D => B, CK => clk, Q => n10, QN => n14
                           );
   MY_CLK_r_REG313_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => n15
                           );
   U1 : XNOR2_X1 port map( A => n14, B => n15, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_399;

architecture SYN_BEHAVIORAL of FA_399 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n10, n11, n12, n14, n15, n16 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n10, B => n6, ZN => S);
   U3 : XNOR2_X1 port map( A => n11, B => n12, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => n5);
   U8 : AOI22_X1 port map( A1 => n5, A2 => n14, B1 => n16, B2 => n15, ZN => Co)
                           ;
   MY_CLK_r_REG175_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n16
                           );
   MY_CLK_r_REG314_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n15
                           );
   MY_CLK_r_REG330_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_400;

architecture SYN_BEHAVIORAL of FA_400 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n5, n8, n9, n11, n12 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => n9, B => n8, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => n9, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n11, B1 => n12, B2 => n1, ZN => Co);
   MY_CLK_r_REG149_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG346_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n11
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_401;

architecture SYN_BEHAVIORAL of FA_401 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n5, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U4 : NAND2_X1 port map( A1 => B, A2 => n10, ZN => n5);
   U7 : INV_X1 port map( A => B, ZN => n2);
   U8 : AOI22_X1 port map( A1 => n5, A2 => n13, B1 => n12, B2 => n2, ZN => Co);
   MY_CLK_r_REG162_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG355_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => n13
                           );
   U1 : XNOR2_X1 port map( A => n9, B => n10, ZN => n14);
   U2 : XNOR2_X1 port map( A => B, B => n14, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_402;

architecture SYN_BEHAVIORAL of FA_402 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n8, n9, n11, n12 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => n9, B => n8, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n11, B1 => n2, B2 => n12, ZN => Co);
   MY_CLK_r_REG356_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG367_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n11
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_403;

architecture SYN_BEHAVIORAL of FA_403 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n9, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n13, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG147_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG368_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG375_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n14
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_404;

architecture SYN_BEHAVIORAL of FA_404 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n8, n9, n10, n_1703, n_1704, n_1705 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => n2);
   U4 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n3);
   U5 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U6 : XNOR2_X1 port map( A => n8, B => n9, ZN => n4);
   MY_CLK_r_REG268_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => 
                           n_1703);
   MY_CLK_r_REG376_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => 
                           n_1704);
   MY_CLK_r_REG364_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1705);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_405;

architecture SYN_BEHAVIORAL of FA_405 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5, n10, n11, n12, n13, n15, n_1706, n_1707, n_1708 : 
      std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n12, B => n11, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n15, B2 => n13, A => n10, ZN => Co);
   MY_CLK_r_REG366_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n13, QN => 
                           n_1706);
   MY_CLK_r_REG280_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n15
                           );
   MY_CLK_r_REG365_S1 : DFF_X1 port map( D => n5, CK => clk, Q => n11, QN => 
                           n_1707);
   MY_CLK_r_REG281_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1708);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_406;

architecture SYN_BEHAVIORAL of FA_406 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n14, A => n1, ZN => Co);
   MY_CLK_r_REG287_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG387_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG362_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_407;

architecture SYN_BEHAVIORAL of FA_407 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1709, n_1710 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG363_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1709);
   MY_CLK_r_REG325_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1710);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_408;

architecture SYN_BEHAVIORAL of FA_408 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6, n7, n_1711, n_1712 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   MY_CLK_r_REG386_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => 
                           n_1711);
   MY_CLK_r_REG294_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n6, QN => 
                           n_1712);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_409;

architecture SYN_BEHAVIORAL of FA_409 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_411;

architecture SYN_BEHAVIORAL of FA_411 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n3, B2 => n4, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_412;

architecture SYN_BEHAVIORAL of FA_412 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n9, n10, n11, n_1713, n_1714, n_1715 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   MY_CLK_r_REG337_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n11, QN => 
                           n_1713);
   MY_CLK_r_REG385_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n10, QN => 
                           n_1714);
   MY_CLK_r_REG338_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n9, QN => 
                           n_1715);
   U1 : OAI21_X1 port map( B1 => n11, B2 => n10, A => n9, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_414;

architecture SYN_BEHAVIORAL of FA_414 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_429;

architecture SYN_BEHAVIORAL of FA_429 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n6, n_1717, n_1718 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n5, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   MY_CLK_r_REG16_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1717);
   MY_CLK_r_REG481_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n5, QN => 
                           n_1718);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_430;

architecture SYN_BEHAVIORAL of FA_430 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_431;

architecture SYN_BEHAVIORAL of FA_431 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_432;

architecture SYN_BEHAVIORAL of FA_432 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5, n10, n11, n12, n13, n15, n_1719, n_1720, n_1721 : 
      std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n11, B => n10, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n10, A2 => n15, B1 => n13, B2 => n12, ZN => Co
                           );
   MY_CLK_r_REG486_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n13, QN => 
                           n_1719);
   MY_CLK_r_REG490_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n12, QN => 
                           n_1720);
   MY_CLK_r_REG225_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n11, QN => 
                           n15);
   MY_CLK_r_REG487_S1 : DFF_X1 port map( D => n5, CK => clk, Q => n10, QN => 
                           n_1721);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_433;

architecture SYN_BEHAVIORAL of FA_433 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6, n7, n_1722, n_1723 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   MY_CLK_r_REG488_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => 
                           n_1722);
   MY_CLK_r_REG480_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n6, QN => 
                           n_1723);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_434;

architecture SYN_BEHAVIORAL of FA_434 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n_1724, n_1725, n_1726 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n3);
   U5 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n2);
   MY_CLK_r_REG489_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1724);
   MY_CLK_r_REG484_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1725);
   MY_CLK_r_REG220_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1726);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_435;

architecture SYN_BEHAVIORAL of FA_435 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n14, A => n1, ZN => Co);
   MY_CLK_r_REG485_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG482_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG222_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_436;

architecture SYN_BEHAVIORAL of FA_436 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n1, ZN => Co);
   MY_CLK_r_REG483_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG212_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG211_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n14
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_437;

architecture SYN_BEHAVIORAL of FA_437 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net30807, n1, n5, n6, n7, n9, n10, n_1727 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n6, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => n5, ZN => S);
   U4 : OAI21_X1 port map( B1 => n6, B2 => n7, A => n5, ZN => net30807);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n9, A => net30807, ZN => Co);
   MY_CLK_r_REG213_S1 : DFF_X1 port map( D => A, CK => clk, Q => n7, QN => n10)
                           ;
   MY_CLK_r_REG202_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => n9);
   MY_CLK_r_REG201_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n5, QN => 
                           n_1727);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_438;

architecture SYN_BEHAVIORAL of FA_438 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n9, n10, n11, n13, n14, n17, n_1728 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => n5);
   U6 : AOI22_X1 port map( A1 => n5, A2 => n13, B1 => n14, B2 => n17, ZN => Co)
                           ;
   U7 : FA_X1 port map( A => n11, B => n10, CI => n9, CO => n_1728, S => S);
   MY_CLK_r_REG203_S1 : DFF_X1 port map( D => A, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG206_S1 : DFF_X1 port map( D => B, CK => clk, Q => n10, QN => n17
                           );
   MY_CLK_r_REG205_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => n13
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_439;

architecture SYN_BEHAVIORAL of FA_439 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n8, B => n7, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n10, B2 => n11, ZN => Co);
   MY_CLK_r_REG207_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG191_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n11)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_440;

architecture SYN_BEHAVIORAL of FA_440 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n8, n9, n10, n12, n13, n_1729 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n2, B => n8, ZN => S);
   U4 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => Co);
   U5 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n4);
   MY_CLK_r_REG190_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG491_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG193_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1729);
   U1 : XNOR2_X1 port map( A => n12, B => n13, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_441;

architecture SYN_BEHAVIORAL of FA_441 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n_1730, n_1731, n_1732 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n1);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n2);
   MY_CLK_r_REG492_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1730);
   MY_CLK_r_REG173_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1731);
   MY_CLK_r_REG172_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1732);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_442;

architecture SYN_BEHAVIORAL of FA_442 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7, n11, n13, n14, n_1733 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => A, B => n7, ZN => S);
   U5 : NAND2_X1 port map( A1 => n11, A2 => A, ZN => n6);
   U7 : INV_X1 port map( A => A, ZN => n4);
   MY_CLK_r_REG177_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG176_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n_1733, QN =>
                           n13);
   U1 : AOI22_X1 port map( A1 => n6, A2 => n13, B1 => n4, B2 => n14, ZN => Co);
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_443;

architecture SYN_BEHAVIORAL of FA_443 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net30829, n2, n6, n7, n8, n10, n11, n12 : std_logic;

begin
   
   U4 : XNOR2_X1 port map( A => n2, B => n6, ZN => S);
   U6 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => net30829);
   MY_CLK_r_REG178_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n11)
                           ;
   MY_CLK_r_REG158_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n12)
                           ;
   MY_CLK_r_REG157_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n10
                           );
   U1 : AOI22_X1 port map( A1 => net30829, A2 => n10, B1 => n11, B2 => n12, ZN 
                           => Co);
   U2 : XNOR2_X1 port map( A => n11, B => n12, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_444;

architecture SYN_BEHAVIORAL of FA_444 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n6, n10, n11, n12, n14, n15, n16 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => n10, ZN => S);
   U7 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => n3);
   MY_CLK_r_REG159_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n15
                           );
   MY_CLK_r_REG161_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n16
                           );
   MY_CLK_r_REG163_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n14);
   U1 : AOI22_X1 port map( A1 => n15, A2 => n16, B1 => n3, B2 => n14, ZN => Co)
                           ;
   U2 : XNOR2_X1 port map( A => n15, B => n16, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_445;

architecture SYN_BEHAVIORAL of FA_445 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n6, n10, n11, n12, n14, n15, n16 : std_logic;

begin
   
   U4 : XNOR2_X1 port map( A => n6, B => n11, ZN => S);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n12, A => n10, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n15, B2 => n14, A => n3, ZN => Co);
   MY_CLK_r_REG160_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n15
                           );
   MY_CLK_r_REG145_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG139_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n16);
   U1 : XNOR2_X1 port map( A => n15, B => n16, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_446;

architecture SYN_BEHAVIORAL of FA_446 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n9, n10, n11, n13, n14, n15 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => n9, ZN => S);
   U4 : NAND2_X1 port map( A1 => n11, A2 => n10, ZN => n4);
   MY_CLK_r_REG146_S1 : DFF_X1 port map( D => A, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG127_S1 : DFF_X1 port map( D => B, CK => clk, Q => n10, QN => n15
                           );
   MY_CLK_r_REG148_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => n13
                           );
   U1 : AOI22_X1 port map( A1 => n4, A2 => n13, B1 => n14, B2 => n15, ZN => Co)
                           ;
   U3 : XNOR2_X1 port map( A => n14, B => n15, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_447;

architecture SYN_BEHAVIORAL of FA_447 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n6, n10, n11, n12, n14, n15, n16 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => n11, ZN => S);
   U7 : OAI21_X1 port map( B1 => n11, B2 => n12, A => n10, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n15, B2 => n14, A => n3, ZN => Co);
   MY_CLK_r_REG136_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n15
                           );
   MY_CLK_r_REG137_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG269_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n16);
   U1 : XNOR2_X1 port map( A => n15, B => n16, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_448;

architecture SYN_BEHAVIORAL of FA_448 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n6, n13, n14, n16, n17, n18, n19, n_1734 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n16, A2 => n18, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n6, A2 => n17, ZN => n2);
   U9 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => n6);
   MY_CLK_r_REG138_S1 : DFF_X1 port map( D => A, CK => clk, Q => n14, QN => n16
                           );
   MY_CLK_r_REG117_S1 : DFF_X1 port map( D => B, CK => clk, Q => n13, QN => n18
                           );
   MY_CLK_r_REG282_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n_1734, QN =>
                           n17);
   U3 : AND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);
   U4 : XNOR2_X1 port map( A => n17, B => n18, ZN => n19);
   U5 : XNOR2_X1 port map( A => n14, B => n19, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_449;

architecture SYN_BEHAVIORAL of FA_449 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n11, n12, n13, n15, n16, n17 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n11, A2 => n16, ZN => n4);
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U3 : XNOR2_X1 port map( A => n4, B => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n11, A2 => n15, ZN => n3);
   U5 : NAND2_X1 port map( A1 => n13, A2 => n12, ZN => n5);
   U7 : XNOR2_X1 port map( A => n7, B => n12, ZN => S);
   MY_CLK_r_REG124_S1 : DFF_X1 port map( D => A, CK => clk, Q => n13, QN => n16
                           );
   MY_CLK_r_REG125_S1 : DFF_X1 port map( D => B, CK => clk, Q => n12, QN => n15
                           );
   MY_CLK_r_REG288_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n11, QN => 
                           n17);
   U8 : XNOR2_X1 port map( A => n16, B => n17, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_450;

architecture SYN_BEHAVIORAL of FA_450 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5, n6, n7, n8, n9, n14, n15, n16, n17, n19, n20, n_1735, n_1736 
      : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n15, B => n14, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => n7, ZN => n9);
   U7 : NAND2_X1 port map( A1 => n17, A2 => n16, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n17, A2 => n20, ZN => n7);
   U9 : NAND2_X1 port map( A1 => n15, A2 => n19, ZN => n8);
   U11 : INV_X1 port map( A => B, ZN => n5);
   MY_CLK_r_REG326_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n17, QN => 
                           n_1735);
   MY_CLK_r_REG103_S1 : DFF_X1 port map( D => n5, CK => clk, Q => n16, QN => 
                           n19);
   MY_CLK_r_REG126_S1 : DFF_X1 port map( D => A, CK => clk, Q => n15, QN => n20
                           );
   MY_CLK_r_REG107_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n14, QN => 
                           n_1736);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_451;

architecture SYN_BEHAVIORAL of FA_451 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n6, n7, n13, n14, n15, n17, n18, n19, n_1737, n_1738 : std_logic;

begin
   
   U5 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);
   U6 : NAND2_X1 port map( A1 => n13, A2 => n15, ZN => n7);
   U7 : INV_X1 port map( A => Ci, ZN => n6);
   MY_CLK_r_REG109_S1 : DFF_X1 port map( D => A, CK => clk, Q => n15, QN => n17
                           );
   MY_CLK_r_REG295_S1 : DFF_X1 port map( D => n6, CK => clk, Q => n14, QN => 
                           n_1737);
   MY_CLK_r_REG81_S1 : DFF_X1 port map( D => B, CK => clk, Q => n13, QN => n19)
                           ;
   MY_CLK_r_REG108_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n_1738, QN =>
                           n18);
   U1 : AOI22_X1 port map( A1 => n14, A2 => n7, B1 => n17, B2 => n19, ZN => Co)
                           ;
   U2 : XNOR2_X1 port map( A => n18, B => n19, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_452;

architecture SYN_BEHAVIORAL of FA_452 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_453;

architecture SYN_BEHAVIORAL of FA_453 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_454;

architecture SYN_BEHAVIORAL of FA_454 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U3 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U4 : INV_X1 port map( A => Ci, ZN => n2);
   U5 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_455;

architecture SYN_BEHAVIORAL of FA_455 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => A, ZN => n3);
   U7 : INV_X1 port map( A => B, ZN => n2);
   U8 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_456;

architecture SYN_BEHAVIORAL of FA_456 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n10, n11, n_1739, n_1740 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG289_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1739, QN => 
                           n10);
   MY_CLK_r_REG297_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n_1740, QN =>
                           n11);
   U2 : XNOR2_X1 port map( A => n10, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_457;

architecture SYN_BEHAVIORAL of FA_457 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n10, n11, n_1741, n_1742 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG305_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1741, QN => 
                           n10);
   MY_CLK_r_REG299_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n_1742, QN =>
                           n11);
   U1 : XNOR2_X1 port map( A => n10, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_458;

architecture SYN_BEHAVIORAL of FA_458 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_460;

architecture SYN_BEHAVIORAL of FA_460 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => B, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_462;

architecture SYN_BEHAVIORAL of FA_462 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_21 is

   port( B : in std_logic;  C, S_BAR : out std_logic;  A_BAR : in std_logic);

end HA_21;

architecture SYN_rtl of HA_21 is

begin
   S_BAR <= A_BAR;

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_465 is

   port( A, B, Ci : in std_logic;  Co : out std_logic;  clk : in std_logic;  
         S_BAR : out std_logic);

end FA_465;

architecture SYN_BEHAVIORAL of FA_465 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n_1748 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   MY_CLK_r_REG315_S1 : DFF_X1 port map( D => n2, CK => clk, Q => S_BAR, QN => 
                           n_1748);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_466 is

   port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_466;

architecture SYN_BEHAVIORAL of FA_466 is

begin
   S_BAR <= A_BAR;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_476 is

   port( Ci : in std_logic;  Co : out std_logic;  B_BAR, A_BAR : in std_logic; 
         S_BAR : out std_logic);

end FA_476;

architecture SYN_BEHAVIORAL of FA_476 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n8, B => A_BAR, Z => S_BAR);
   U1 : NOR2_X1 port map( A1 => A_BAR, A2 => B_BAR, ZN => Co);
   U3 : INV_X1 port map( A => B_BAR, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_478 is

   port( A, B, Ci : in std_logic;  S : out std_logic;  clk : in std_logic;  
         Co_BAR : out std_logic);

end FA_478;

architecture SYN_BEHAVIORAL of FA_478 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n6, n_1754, n_1755 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n3, A2 => n6, ZN => Co_BAR);
   U5 : XOR2_X1 port map( A => n6, B => n3, Z => S);
   MY_CLK_r_REG449_S1 : DFF_X1 port map( D => A, CK => clk, Q => n3, QN => 
                           n_1754);
   MY_CLK_r_REG459_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => 
                           n_1755);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_479 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_479;

architecture SYN_BEHAVIORAL of FA_479 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_482 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_482;

architecture SYN_BEHAVIORAL of FA_482 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_483;

architecture SYN_BEHAVIORAL of FA_483 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_22 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_22;

architecture SYN_rtl of HA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_486 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_486;

architecture SYN_BEHAVIORAL of FA_486 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_490 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_490;

architecture SYN_BEHAVIORAL of FA_490 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_491 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_491;

architecture SYN_BEHAVIORAL of FA_491 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_492 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_492;

architecture SYN_BEHAVIORAL of FA_492 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_493 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_493;

architecture SYN_BEHAVIORAL of FA_493 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_494;

architecture SYN_BEHAVIORAL of FA_494 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U5 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_495;

architecture SYN_BEHAVIORAL of FA_495 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_496;

architecture SYN_BEHAVIORAL of FA_496 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1756, n_1757 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG345_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1756);
   MY_CLK_r_REG331_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1757);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_497;

architecture SYN_BEHAVIORAL of FA_497 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1758, n_1759 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG354_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1758);
   MY_CLK_r_REG347_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1759);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_498;

architecture SYN_BEHAVIORAL of FA_498 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_499;

architecture SYN_BEHAVIORAL of FA_499 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_500;

architecture SYN_BEHAVIORAL of FA_500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n2, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : AOI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U7 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_501;

architecture SYN_BEHAVIORAL of FA_501 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_506;

architecture SYN_BEHAVIORAL of FA_506 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n2, B2 => n3, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_508;

architecture SYN_BEHAVIORAL of FA_508 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_509;

architecture SYN_BEHAVIORAL of FA_509 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_510;

architecture SYN_BEHAVIORAL of FA_510 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_511;

architecture SYN_BEHAVIORAL of FA_511 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_518 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_518;

architecture SYN_BEHAVIORAL of FA_518 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_519 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_519;

architecture SYN_BEHAVIORAL of FA_519 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n10, n11, n_1761, n_1762 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG270_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n_1761, QN =>
                           n10);
   MY_CLK_r_REG189_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n_1762, QN =>
                           n11);
   U1 : XNOR2_X1 port map( A => n10, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_520 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_520;

architecture SYN_BEHAVIORAL of FA_520 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n2, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n2);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U1 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_521 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_521;

architecture SYN_BEHAVIORAL of FA_521 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : AOI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_522 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_522;

architecture SYN_BEHAVIORAL of FA_522 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_523 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_523;

architecture SYN_BEHAVIORAL of FA_523 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_524 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_524;

architecture SYN_BEHAVIORAL of FA_524 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_525 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_525;

architecture SYN_BEHAVIORAL of FA_525 is

   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n17, n_1763, n_1764, 
      n_1765 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n9, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => A, ZN => n9);
   U5 : INV_X1 port map( A => A, ZN => n8);
   U6 : INV_X1 port map( A => B, ZN => n7);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U8 : INV_X1 port map( A => Ci, ZN => n3);
   U9 : NOR2_X1 port map( A1 => A, A2 => n3, ZN => n4);
   U10 : XOR2_X1 port map( A => n5, B => n4, Z => n6);
   U11 : OAI21_X1 port map( B1 => n15, B2 => n14, A => n13, ZN => Co);
   MY_CLK_r_REG143_S1 : DFF_X1 port map( D => n8, CK => clk, Q => n15, QN => 
                           n_1763);
   MY_CLK_r_REG144_S1 : DFF_X1 port map( D => n6, CK => clk, Q => n13, QN => 
                           n_1764);
   MY_CLK_r_REG302_S1 : SDFF_X1 port map( D => n7, SI => n17, SE => n17, CK => 
                           clk, Q => n14, QN => n_1765);
   n17 <= '0';

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_526 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_526;

architecture SYN_BEHAVIORAL of FA_526 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n7 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => A, B => n7, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_527 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_527;

architecture SYN_BEHAVIORAL of FA_527 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_528 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_528;

architecture SYN_BEHAVIORAL of FA_528 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_529 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_529;

architecture SYN_BEHAVIORAL of FA_529 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_534 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_534;

architecture SYN_BEHAVIORAL of FA_534 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_535 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_535;

architecture SYN_BEHAVIORAL of FA_535 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_536 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_536;

architecture SYN_BEHAVIORAL of FA_536 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_539 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic);

end FA_539;

architecture SYN_BEHAVIORAL of FA_539 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => A_BAR, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_541 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic);

end FA_541;

architecture SYN_BEHAVIORAL of FA_541 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n6, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => A_BAR, B2 => n1, ZN => Co)
                           ;
   U3 : INV_X1 port map( A => A_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_543 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic);

end FA_543;

architecture SYN_BEHAVIORAL of FA_543 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => n6, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => B_BAR, ZN => Co)
                           ;
   U5 : INV_X1 port map( A => B_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_544 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_544;

architecture SYN_BEHAVIORAL of FA_544 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_546 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_546;

architecture SYN_BEHAVIORAL of FA_546 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_547 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_547;

architecture SYN_BEHAVIORAL of FA_547 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net31297, net31298, net31299, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net31299);
   U4 : INV_X1 port map( A => A, ZN => net31297);
   U5 : INV_X1 port map( A => B, ZN => net31298);
   U6 : OAI21_X1 port map( B1 => net31297, B2 => net31298, A => net31299, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_549 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_549;

architecture SYN_BEHAVIORAL of FA_549 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n1);
   U2 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_550 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_550;

architecture SYN_BEHAVIORAL of FA_550 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_551 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_551;

architecture SYN_BEHAVIORAL of FA_551 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_552 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_552;

architecture SYN_BEHAVIORAL of FA_552 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n10, n11, n_1767, n_1768 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG495_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1767, QN => 
                           n10);
   MY_CLK_r_REG174_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n_1768, QN =>
                           n11);
   U1 : XNOR2_X1 port map( A => n10, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_553 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_553;

architecture SYN_BEHAVIORAL of FA_553 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net31320, net31321, net31322, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net31322);
   U4 : INV_X1 port map( A => B, ZN => net31321);
   U5 : INV_X1 port map( A => A, ZN => net31320);
   U7 : OAI21_X1 port map( B1 => net31320, B2 => net31321, A => net31322, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_554 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_554;

architecture SYN_BEHAVIORAL of FA_554 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_555 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_555;

architecture SYN_BEHAVIORAL of FA_555 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n6, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n6);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : INV_X1 port map( A => B, ZN => n4);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U7 : INV_X1 port map( A => Ci, ZN => n2);
   U8 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_556 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_556;

architecture SYN_BEHAVIORAL of FA_556 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_557 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_557;

architecture SYN_BEHAVIORAL of FA_557 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => A, ZN => n4);
   U8 : INV_X1 port map( A => B, ZN => n3);
   U9 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_558 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_558;

architecture SYN_BEHAVIORAL of FA_558 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U7 : INV_X1 port map( A => Ci, ZN => n1);
   U1 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_559 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_559;

architecture SYN_BEHAVIORAL of FA_559 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_560 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_560;

architecture SYN_BEHAVIORAL of FA_560 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_562 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_562;

architecture SYN_BEHAVIORAL of FA_562 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n7 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => n7, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_563 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_563;

architecture SYN_BEHAVIORAL of FA_563 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_565 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_565;

architecture SYN_BEHAVIORAL of FA_565 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_566 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_566;

architecture SYN_BEHAVIORAL of FA_566 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : INV_X1 port map( A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U5 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_567 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_567;

architecture SYN_BEHAVIORAL of FA_567 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_33 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_33;

architecture SYN_rtl of HA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);
   U2 : XOR2_X1 port map( A => A, B => B, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_569 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_569;

architecture SYN_BEHAVIORAL of FA_569 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_570 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_570;

architecture SYN_BEHAVIORAL of FA_570 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_571 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_571;

architecture SYN_BEHAVIORAL of FA_571 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_572 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_572;

architecture SYN_BEHAVIORAL of FA_572 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_573 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_573;

architecture SYN_BEHAVIORAL of FA_573 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_574 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_574;

architecture SYN_BEHAVIORAL of FA_574 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_576 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_576;

architecture SYN_BEHAVIORAL of FA_576 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_577 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_577;

architecture SYN_BEHAVIORAL of FA_577 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n1);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U3 : OAI22_X1 port map( A1 => n2, A2 => n1, B1 => Ci, B2 => n2, ZN => n3);
   U4 : INV_X1 port map( A => n3, ZN => Co);
   U5 : XOR2_X1 port map( A => Ci, B => n1, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_578 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_578;

architecture SYN_BEHAVIORAL of FA_578 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U5 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_579 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_579;

architecture SYN_BEHAVIORAL of FA_579 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_580 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_580;

architecture SYN_BEHAVIORAL of FA_580 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U2 : OR2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n1, A2 => Ci, ZN => n4);
   U4 : XNOR2_X1 port map( A => n2, B => Ci, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n2);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_581 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_581;

architecture SYN_BEHAVIORAL of FA_581 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_582 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_582;

architecture SYN_BEHAVIORAL of FA_582 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_583 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_583;

architecture SYN_BEHAVIORAL of FA_583 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_584 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_584;

architecture SYN_BEHAVIORAL of FA_584 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_585 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_585;

architecture SYN_BEHAVIORAL of FA_585 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_587 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_587;

architecture SYN_BEHAVIORAL of FA_587 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_588 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_588;

architecture SYN_BEHAVIORAL of FA_588 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_589 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_589;

architecture SYN_BEHAVIORAL of FA_589 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => A, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => B, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_590 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_590;

architecture SYN_BEHAVIORAL of FA_590 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U2 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n1);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_591 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_591;

architecture SYN_BEHAVIORAL of FA_591 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => B, ZN => n3);
   U4 : INV_X1 port map( A => A, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_592 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_592;

architecture SYN_BEHAVIORAL of FA_592 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U2 : XOR2_X1 port map( A => A, B => n1, Z => S);
   U3 : XOR2_X1 port map( A => B, B => Ci, Z => n1);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_42 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_42;

architecture SYN_rtl of HA_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   C <= B;
   
   U1 : INV_X1 port map( A => B, ZN => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_593 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_593;

architecture SYN_BEHAVIORAL of FA_593 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : AOI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_594 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_594;

architecture SYN_BEHAVIORAL of FA_594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_595 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_595;

architecture SYN_BEHAVIORAL of FA_595 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net31526, net31527, net31528, net31529, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U3 : INV_X1 port map( A => B, ZN => net31529);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net31526);
   U5 : INV_X1 port map( A => Ci, ZN => net31527);
   U6 : INV_X1 port map( A => A, ZN => net31528);
   U7 : AOI22_X1 port map( A1 => net31526, A2 => net31527, B1 => net31528, B2 
                           => net31529, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_596 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_596;

architecture SYN_BEHAVIORAL of FA_596 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => B, B2 => n3, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_597 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_597;

architecture SYN_BEHAVIORAL of FA_597 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_598 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_598;

architecture SYN_BEHAVIORAL of FA_598 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n6 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => S);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n6, A => Ci, ZN => n2);
   U1 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   n6 <= '1';

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_599 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic);

end FA_599;

architecture SYN_BEHAVIORAL of FA_599 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => n6, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => B_BAR, ZN => Co)
                           ;
   U5 : INV_X1 port map( A => B_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_600 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic);

end FA_600;

architecture SYN_BEHAVIORAL of FA_600 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => A_BAR, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => A_BAR, B2 => n1, ZN => Co)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_601 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_601;

architecture SYN_BEHAVIORAL of FA_601 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net31554, net31555, net31556, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);
   U3 : INV_X1 port map( A => B, ZN => net31555);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net31556);
   U5 : INV_X1 port map( A => A, ZN => net31554);
   U6 : OAI21_X1 port map( B1 => net31554, B2 => net31555, A => net31556, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_602 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_602;

architecture SYN_BEHAVIORAL of FA_602 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_603 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_603;

architecture SYN_BEHAVIORAL of FA_603 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_604 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_604;

architecture SYN_BEHAVIORAL of FA_604 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U5 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_605 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_605;

architecture SYN_BEHAVIORAL of FA_605 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U3 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_606 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_606;

architecture SYN_BEHAVIORAL of FA_606 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U5 : AOI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_607 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_607;

architecture SYN_BEHAVIORAL of FA_607 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U2 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_43 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_43;

architecture SYN_rtl of HA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_0 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_0;

architecture SYN_rtl of HA_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_1 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
         p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
         p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
         p_17_port, p_16_port, p_15_port, p_14_BAR, p_13_port, p_12_port, 
         p_11_port, p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, p_5_port
         , p_4_port, p_3_port, p_2_port, p_1_port, p_0_port : out std_logic);

end ENC_1;

architecture SYN_beh of ENC_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n56, n58, n59, n68, n69, n85, n118, n120, n134, n_1837 : std_logic;

begin
   
   U87 : MUX2_X1 port map( A => n69, B => n134, S => A(14), Z => n56);
   U89 : MUX2_X1 port map( A => n118, B => n85, S => A(14), Z => n59);
   U90 : MUX2_X1 port map( A => n68, B => n120, S => A(15), Z => n58);
   MY_CLK_r_REG351_S1 : DFF_X1 port map( D => n56, CK => clk, Q => p_14_BAR, QN
                           => n_1837);
   n68 <= '1';
   n69 <= '1';
   n85 <= '1';
   n118 <= '1';
   n120 <= '1';
   n134 <= '1';
   U3 : NAND2_X1 port map( A1 => n59, A2 => n58, ZN => p_15_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_2 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
         p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
         p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
         p_17_port, p_16_BAR, p_15_port, p_14_port, p_13_port, p_12_port, 
         p_11_port, p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, p_5_port
         , p_4_port, p_3_port, p_2_port, p_1_port, p_0_port : out std_logic);

end ENC_2;

architecture SYN_beh of ENC_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n60, n62, n63, n75, n76, n99, n131, n134, n135, n_1902 : std_logic;

begin
   
   U91 : MUX2_X1 port map( A => n76, B => n134, S => A(16), Z => n60);
   U93 : MUX2_X1 port map( A => n131, B => n99, S => A(16), Z => n63);
   U94 : MUX2_X1 port map( A => n75, B => n135, S => A(17), Z => n62);
   MY_CLK_r_REG336_S1 : DFF_X1 port map( D => n60, CK => clk, Q => p_16_BAR, QN
                           => n_1902);
   n75 <= '1';
   n76 <= '1';
   n99 <= '1';
   n131 <= '1';
   n134 <= '1';
   n135 <= '1';
   U3 : NAND2_X1 port map( A1 => n63, A2 => n62, ZN => p_17_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_3 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
         p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
         p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
         p_17_port, p_15_port, p_14_port, p_13_port, p_12_port, p_11_port, 
         p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, p_5_port, p_4_BAR, 
         p_3_port, p_2_port, p_1_port, p_0_port, p_16_BAR : out std_logic);

end ENC_3;

architecture SYN_beh of ENC_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n24, n27, n28, n30, n31, n32, n33, n35, n59, n61, n62, n63, n64, n65,
      n66, n16, n17, n18, n19, n86, n87, n88, n98, n107, n108, n109, n116, n117
      , n118, n119, n120, n121, n122, n123, n130, n131, n132, n145, n146, n147,
      n148, n161, n162, n163, n164, n_1954, n_1955 : std_logic;

begin
   
   U36 : MUX2_X1 port map( A => n148, B => n119, S => A(0), Z => n24);
   U39 : MUX2_X1 port map( A => n86, B => n164, S => A(0), Z => n28);
   U42 : MUX2_X1 port map( A => n163, B => n118, S => A(1), Z => n27);
   U44 : MUX2_X1 port map( A => n98, B => n147, S => A(1), Z => n31);
   U46 : MUX2_X1 port map( A => n162, B => n117, S => A(2), Z => n30);
   U48 : MUX2_X1 port map( A => n87, B => n146, S => A(2), Z => n33);
   U49 : MUX2_X1 port map( A => n161, B => n116, S => A(3), Z => n32);
   U51 : MUX2_X1 port map( A => n88, B => n145, S => A(3), Z => n35);
   U88 : MUX2_X1 port map( A => n19, B => n123, S => A(16), Z => n59);
   U90 : MUX2_X1 port map( A => n107, B => n132, S => A(16), Z => n62);
   U91 : MUX2_X1 port map( A => n18, B => n122, S => A(17), Z => n61);
   U93 : MUX2_X1 port map( A => n108, B => n131, S => A(17), Z => n64);
   U94 : MUX2_X1 port map( A => n17, B => n121, S => A(18), Z => n63);
   U96 : MUX2_X1 port map( A => n109, B => n130, S => A(18), Z => n66);
   U97 : MUX2_X1 port map( A => n16, B => n120, S => A(19), Z => n65);
   MY_CLK_r_REG453_S1 : DFF_X1 port map( D => n35, CK => clk, Q => p_4_BAR, QN 
                           => n_1954);
   MY_CLK_r_REG335_S1 : DFF_X1 port map( D => n59, CK => clk, Q => p_16_BAR, QN
                           => n_1955);
   n16 <= '1';
   n17 <= '1';
   n18 <= '1';
   n19 <= '1';
   n86 <= '1';
   n87 <= '1';
   n88 <= '1';
   n98 <= '1';
   n107 <= '1';
   n108 <= '1';
   n109 <= '1';
   n116 <= '1';
   n117 <= '1';
   n118 <= '1';
   n119 <= '1';
   n120 <= '1';
   n121 <= '1';
   n122 <= '1';
   n123 <= '1';
   n130 <= '1';
   n131 <= '1';
   n132 <= '1';
   n145 <= '1';
   n146 <= '1';
   n147 <= '1';
   n148 <= '1';
   n161 <= '1';
   n162 <= '1';
   n163 <= '1';
   n164 <= '1';
   U7 : NAND2_X1 port map( A1 => n31, A2 => n30, ZN => p_2_port);
   U8 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => p_17_port);
   U9 : NAND2_X1 port map( A1 => n33, A2 => n32, ZN => p_3_port);
   U10 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => p_18_port);
   U11 : NAND2_X1 port map( A1 => n28, A2 => n27, ZN => p_1_port);
   U12 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => p_19_port);
   U13 : INV_X1 port map( A => n24, ZN => p_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_4 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
         p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
         p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
         p_17_port, p_15_port, p_14_port, p_13_port, p_12_port, p_11_port, 
         p_10_port, p_9_port, p_8_port, p_7_port, p_6_BAR, p_5_port, p_4_port, 
         p_3_port, p_2_port, p_1_port, p_0_port, p_16_BAR : out std_logic);

end ENC_4;

architecture SYN_beh of ENC_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n26, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n40, n60, n61,
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n88, n90, n92, n96, n97, n98
      , n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n120,
      n121, n123, n124, n125, n126, n127, n130, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n162, n164, n165, n176, 
      n177, n178, n179, n180, n_1999, n_2000 : std_logic;

begin
   
   U36 : MUX2_X1 port map( A => n121, B => n108, S => A(0), Z => n26);
   U38 : MUX2_X1 port map( A => n123, B => n165, S => A(0), Z => n30);
   U41 : MUX2_X1 port map( A => n180, B => n107, S => A(1), Z => n29);
   U43 : MUX2_X1 port map( A => n130, B => n147, S => A(1), Z => n32);
   U44 : MUX2_X1 port map( A => n179, B => n106, S => A(2), Z => n31);
   U46 : MUX2_X1 port map( A => n124, B => n148, S => A(2), Z => n34);
   U47 : MUX2_X1 port map( A => n178, B => n105, S => A(3), Z => n33);
   U49 : MUX2_X1 port map( A => n125, B => n149, S => A(3), Z => n36);
   U50 : MUX2_X1 port map( A => n177, B => n104, S => A(4), Z => n35);
   U52 : MUX2_X1 port map( A => n126, B => n150, S => A(4), Z => n38);
   U53 : MUX2_X1 port map( A => n176, B => n103, S => A(5), Z => n37);
   U55 : MUX2_X1 port map( A => n127, B => n151, S => A(5), Z => n40);
   U85 : MUX2_X1 port map( A => n98, B => n113, S => A(16), Z => n60);
   U88 : MUX2_X1 port map( A => n139, B => n162, S => A(16), Z => n62);
   U89 : MUX2_X1 port map( A => n97, B => n112, S => A(17), Z => n61);
   U91 : MUX2_X1 port map( A => n140, B => n144, S => A(17), Z => n64);
   U92 : MUX2_X1 port map( A => n96, B => n111, S => A(18), Z => n63);
   U94 : MUX2_X1 port map( A => n141, B => n145, S => A(18), Z => n66);
   U95 : MUX2_X1 port map( A => n92, B => n110, S => A(19), Z => n65);
   U97 : MUX2_X1 port map( A => n142, B => n146, S => A(19), Z => n68);
   U98 : MUX2_X1 port map( A => n90, B => n109, S => A(20), Z => n67);
   U100 : MUX2_X1 port map( A => n143, B => n164, S => A(20), Z => n70);
   U101 : MUX2_X1 port map( A => n88, B => n120, S => A(21), Z => n69);
   MY_CLK_r_REG439_S1 : DFF_X1 port map( D => n40, CK => clk, Q => p_6_BAR, QN 
                           => n_1999);
   MY_CLK_r_REG334_S1 : DFF_X1 port map( D => n60, CK => clk, Q => p_16_BAR, QN
                           => n_2000);
   n88 <= '1';
   n90 <= '1';
   n92 <= '1';
   n96 <= '1';
   n97 <= '1';
   n98 <= '1';
   n103 <= '1';
   n104 <= '1';
   n105 <= '1';
   n106 <= '1';
   n107 <= '1';
   n108 <= '1';
   n109 <= '1';
   n110 <= '1';
   n111 <= '1';
   n112 <= '1';
   n113 <= '1';
   n120 <= '1';
   n121 <= '1';
   n123 <= '1';
   n124 <= '1';
   n125 <= '1';
   n126 <= '1';
   n127 <= '1';
   n130 <= '1';
   n139 <= '1';
   n140 <= '1';
   n141 <= '1';
   n142 <= '1';
   n143 <= '1';
   n144 <= '1';
   n145 <= '1';
   n146 <= '1';
   n147 <= '1';
   n148 <= '1';
   n149 <= '1';
   n150 <= '1';
   n151 <= '1';
   n162 <= '1';
   n164 <= '1';
   n165 <= '1';
   n176 <= '1';
   n177 <= '1';
   n178 <= '1';
   n179 <= '1';
   n180 <= '1';
   U3 : NAND2_X1 port map( A1 => n36, A2 => n35, ZN => p_4_port);
   U4 : NAND2_X1 port map( A1 => n38, A2 => n37, ZN => p_5_port);
   U5 : NAND2_X1 port map( A1 => n32, A2 => n31, ZN => p_2_port);
   U6 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => p_3_port);
   U7 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => p_19_port);
   U8 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => p_18_port);
   U9 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => p_17_port);
   U10 : NAND2_X1 port map( A1 => n30, A2 => n29, ZN => p_1_port);
   U11 : NAND2_X1 port map( A1 => n70, A2 => n69, ZN => p_21_port);
   U12 : NAND2_X1 port map( A1 => n68, A2 => n67, ZN => p_20_port);
   U13 : INV_X1 port map( A => n26, ZN => p_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_5 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_5;

architecture SYN_beh of ENC_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n25, n26, n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n70, n71, n72, n87, n96, n99 : std_logic;

begin
   
   U38 : MUX2_X1 port map( A => n99, B => n99, S => A(0), Z => n26);
   U45 : MUX2_X1 port map( A => n99, B => n99, S => A(1), Z => n28);
   U48 : MUX2_X1 port map( A => n99, B => n99, S => A(2), Z => n31);
   U52 : MUX2_X1 port map( A => n99, B => n99, S => A(3), Z => n33);
   U56 : MUX2_X1 port map( A => n99, B => n99, S => A(4), Z => n34);
   U58 : MUX2_X1 port map( A => n99, B => n99, S => A(5), Z => n37);
   U62 : MUX2_X1 port map( A => n99, B => n99, S => A(6), Z => n39);
   U64 : MUX2_X1 port map( A => n99, B => n99, S => A(7), Z => n42);
   U67 : MUX2_X1 port map( A => n99, B => n99, S => A(8), Z => n44);
   U70 : MUX2_X1 port map( A => n99, B => n99, S => A(9), Z => n46);
   U73 : MUX2_X1 port map( A => n99, B => n99, S => A(10), Z => n48);
   U76 : MUX2_X1 port map( A => n99, B => n99, S => A(11), Z => n50);
   U79 : MUX2_X1 port map( A => n99, B => n99, S => A(12), Z => n52);
   U82 : MUX2_X1 port map( A => n99, B => n99, S => A(13), Z => n54);
   U85 : MUX2_X1 port map( A => n99, B => n99, S => A(14), Z => n56);
   U88 : MUX2_X1 port map( A => n99, B => n99, S => A(15), Z => n58);
   U91 : MUX2_X1 port map( A => n99, B => n99, S => A(16), Z => n60);
   U94 : MUX2_X1 port map( A => n99, B => n99, S => A(17), Z => n62);
   U97 : MUX2_X1 port map( A => n99, B => n99, S => A(18), Z => n64);
   U100 : MUX2_X1 port map( A => n99, B => n99, S => A(19), Z => n66);
   U104 : MUX2_X1 port map( A => n99, B => n99, S => A(20), Z => n67);
   U106 : MUX2_X1 port map( A => n99, B => n99, S => A(21), Z => n70);
   U109 : MUX2_X1 port map( A => n99, B => n99, S => A(22), Z => n72);
   U3 : INV_X1 port map( A => n87, ZN => n2);
   U4 : NAND2_X1 port map( A1 => n33, A2 => n32, ZN => p(4));
   U5 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => p(5));
   U6 : NAND2_X1 port map( A1 => n68, A2 => n67, ZN => p(21));
   U7 : NAND2_X1 port map( A1 => A(7), A2 => n2, ZN => n40);
   U8 : NAND2_X1 port map( A1 => A(1), A2 => n2, ZN => n25);
   U9 : NAND2_X1 port map( A1 => A(3), A2 => n2, ZN => n30);
   U10 : NAND2_X1 port map( A1 => A(21), A2 => n96, ZN => n68);
   U11 : NAND2_X1 port map( A1 => A(4), A2 => n2, ZN => n32);
   U12 : NAND2_X1 port map( A1 => A(5), A2 => n2, ZN => n35);
   U13 : NAND2_X1 port map( A1 => A(22), A2 => n96, ZN => n69);
   U14 : NAND2_X1 port map( A1 => A(20), A2 => n96, ZN => n65);
   U15 : NAND2_X1 port map( A1 => A(8), A2 => n2, ZN => n41);
   U16 : NAND2_X1 port map( A1 => n40, A2 => n39, ZN => p(7));
   U17 : NAND2_X1 port map( A1 => A(2), A2 => n2, ZN => n27);
   U18 : NAND2_X1 port map( A1 => n70, A2 => n69, ZN => p(22));
   U19 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => p(20));
   U20 : NAND2_X1 port map( A1 => n28, A2 => n27, ZN => p(2));
   U21 : NAND2_X1 port map( A1 => n26, A2 => n25, ZN => p(1));
   U22 : AND2_X1 port map( A1 => A(0), A2 => n96, ZN => p(0));
   U24 : INV_X1 port map( A => b(0), ZN => n87);
   U25 : NAND2_X1 port map( A1 => n31, A2 => n30, ZN => p(3));
   U26 : NAND2_X1 port map( A1 => n37, A2 => n36, ZN => p(6));
   U27 : NAND2_X1 port map( A1 => n44, A2 => n43, ZN => p(9));
   U28 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => p(8));
   U29 : NAND2_X1 port map( A1 => n48, A2 => n47, ZN => p(11));
   U30 : NAND2_X1 port map( A1 => n46, A2 => n45, ZN => p(10));
   U31 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => p(12));
   U32 : NAND2_X1 port map( A1 => n52, A2 => n51, ZN => p(13));
   U33 : NAND2_X1 port map( A1 => n54, A2 => n53, ZN => p(14));
   U34 : NAND2_X1 port map( A1 => n56, A2 => n55, ZN => p(15));
   U35 : NAND2_X1 port map( A1 => n58, A2 => n57, ZN => p(16));
   U36 : NAND2_X1 port map( A1 => n60, A2 => n59, ZN => p(17));
   U37 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => p(18));
   U39 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => p(19));
   U40 : NAND2_X1 port map( A1 => n72, A2 => n71, ZN => p(23));
   U41 : NAND2_X1 port map( A1 => A(23), A2 => n96, ZN => n71);
   U42 : INV_X1 port map( A => n87, ZN => n96);
   U43 : NAND2_X1 port map( A1 => A(19), A2 => n2, ZN => n63);
   U44 : NAND2_X1 port map( A1 => A(18), A2 => n96, ZN => n61);
   U47 : NAND2_X1 port map( A1 => A(17), A2 => n96, ZN => n59);
   U49 : NAND2_X1 port map( A1 => A(16), A2 => n96, ZN => n57);
   U50 : NAND2_X1 port map( A1 => A(15), A2 => n96, ZN => n55);
   U51 : NAND2_X1 port map( A1 => A(14), A2 => n96, ZN => n53);
   U53 : NAND2_X1 port map( A1 => A(13), A2 => n96, ZN => n51);
   U54 : NAND2_X1 port map( A1 => A(12), A2 => n2, ZN => n49);
   U55 : NAND2_X1 port map( A1 => A(11), A2 => n2, ZN => n47);
   U57 : NAND2_X1 port map( A1 => A(10), A2 => n2, ZN => n45);
   U59 : NAND2_X1 port map( A1 => A(9), A2 => n2, ZN => n43);
   U60 : NAND2_X1 port map( A1 => A(6), A2 => n2, ZN => n36);
   n99 <= '1';

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_6 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_6;

architecture SYN_beh of ENC_6 is

   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n15, n16, n23, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, 
      n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84, n95, n97, n99, n100, n101, n104, n105 : 
      std_logic;

begin
   
   U3 : AND2_X1 port map( A1 => n62, A2 => n61, ZN => n1);
   U16 : NAND3_X1 port map( A1 => b(0), A2 => n30, A3 => b(1), ZN => n4);
   U20 : NAND2_X1 port map( A1 => n16, A2 => n1, ZN => p(14));
   U33 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n27);
   U37 : INV_X1 port map( A => b(2), ZN => n30);
   U38 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n29);
   U42 : NAND2_X1 port map( A1 => b(2), A2 => n29, ZN => n33);
   U43 : MUX2_X1 port map( A => n33, B => n104, S => A(0), Z => n28);
   U44 : OAI211_X1 port map( C1 => n30, C2 => n29, A => n100, B => n28, ZN => 
                           p(0));
   U45 : NAND3_X1 port map( A1 => n30, A2 => b(0), A3 => b(1), ZN => n101);
   U46 : MUX2_X1 port map( A => n100, B => n23, S => A(0), Z => n36);
   U47 : NAND2_X1 port map( A1 => n32, A2 => n31, ZN => n34);
   U48 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n4, A4 => n95, ZN => 
                           n97);
   U49 : NAND2_X1 port map( A1 => b(2), A2 => n34, ZN => n99);
   U50 : MUX2_X1 port map( A => n99, B => n104, S => A(1), Z => n35);
   U51 : NAND3_X1 port map( A1 => n36, A2 => n97, A3 => n35, ZN => p(1));
   U52 : MUX2_X1 port map( A => n100, B => n23, S => A(1), Z => n38);
   U53 : MUX2_X1 port map( A => n99, B => n104, S => A(2), Z => n37);
   U54 : NAND3_X1 port map( A1 => n38, A2 => n15, A3 => n37, ZN => p(2));
   U55 : MUX2_X1 port map( A => n100, B => n101, S => A(2), Z => n40);
   U56 : MUX2_X1 port map( A => n99, B => n104, S => A(3), Z => n39);
   U57 : NAND3_X1 port map( A1 => n40, A2 => n15, A3 => n39, ZN => p(3));
   U58 : MUX2_X1 port map( A => n100, B => n101, S => A(3), Z => n42);
   U59 : MUX2_X1 port map( A => n99, B => n104, S => A(4), Z => n41);
   U60 : NAND3_X1 port map( A1 => n42, A2 => n97, A3 => n41, ZN => p(4));
   U61 : MUX2_X1 port map( A => n99, B => n95, S => A(5), Z => n44);
   U62 : MUX2_X1 port map( A => n100, B => n23, S => A(4), Z => n43);
   U63 : NAND3_X1 port map( A1 => n44, A2 => n15, A3 => n43, ZN => p(5));
   U64 : MUX2_X1 port map( A => n100, B => n23, S => A(5), Z => n46);
   U65 : MUX2_X1 port map( A => n99, B => n104, S => A(6), Z => n45);
   U66 : NAND3_X1 port map( A1 => n46, A2 => n15, A3 => n45, ZN => p(6));
   U67 : MUX2_X1 port map( A => n100, B => n101, S => A(6), Z => n48);
   U68 : MUX2_X1 port map( A => n99, B => n104, S => A(7), Z => n47);
   U69 : NAND3_X1 port map( A1 => n48, A2 => n15, A3 => n47, ZN => p(7));
   U70 : MUX2_X1 port map( A => n100, B => n101, S => A(7), Z => n50);
   U71 : MUX2_X1 port map( A => n99, B => n95, S => A(8), Z => n49);
   U72 : NAND3_X1 port map( A1 => n50, A2 => n97, A3 => n49, ZN => p(8));
   U73 : MUX2_X1 port map( A => n100, B => n101, S => A(8), Z => n52);
   U74 : MUX2_X1 port map( A => n99, B => n95, S => A(9), Z => n51);
   U75 : NAND3_X1 port map( A1 => n52, A2 => n15, A3 => n51, ZN => p(9));
   U76 : MUX2_X1 port map( A => n100, B => n101, S => A(9), Z => n54);
   U77 : MUX2_X1 port map( A => n99, B => n104, S => A(10), Z => n53);
   U78 : NAND3_X1 port map( A1 => n15, A2 => n54, A3 => n53, ZN => p(10));
   U79 : MUX2_X1 port map( A => n100, B => n101, S => A(10), Z => n56);
   U80 : MUX2_X1 port map( A => n99, B => n104, S => A(11), Z => n55);
   U81 : NAND3_X1 port map( A1 => n56, A2 => n16, A3 => n55, ZN => p(11));
   U82 : MUX2_X1 port map( A => n100, B => n101, S => A(11), Z => n58);
   U83 : MUX2_X1 port map( A => n99, B => n104, S => A(12), Z => n57);
   U84 : NAND3_X1 port map( A1 => n58, A2 => n15, A3 => n57, ZN => p(12));
   U85 : MUX2_X1 port map( A => n100, B => n101, S => A(12), Z => n60);
   U86 : MUX2_X1 port map( A => n99, B => n95, S => A(13), Z => n59);
   U87 : NAND3_X1 port map( A1 => n60, A2 => n16, A3 => n59, ZN => p(13));
   U88 : MUX2_X1 port map( A => n99, B => n104, S => A(14), Z => n62);
   U89 : MUX2_X1 port map( A => n100, B => n4, S => A(13), Z => n61);
   U90 : MUX2_X1 port map( A => n100, B => n23, S => A(14), Z => n64);
   U91 : MUX2_X1 port map( A => n99, B => n104, S => A(15), Z => n63);
   U92 : NAND3_X1 port map( A1 => n64, A2 => n15, A3 => n63, ZN => p(15));
   U93 : MUX2_X1 port map( A => n100, B => n101, S => A(15), Z => n66);
   U94 : MUX2_X1 port map( A => n99, B => n95, S => A(16), Z => n65);
   U95 : NAND3_X1 port map( A1 => n66, A2 => n97, A3 => n65, ZN => p(16));
   U96 : MUX2_X1 port map( A => n100, B => n23, S => A(16), Z => n68);
   U97 : MUX2_X1 port map( A => n99, B => n95, S => A(17), Z => n67);
   U98 : NAND3_X1 port map( A1 => n68, A2 => n15, A3 => n67, ZN => p(17));
   U99 : MUX2_X1 port map( A => n100, B => n23, S => A(17), Z => n70);
   U100 : MUX2_X1 port map( A => n99, B => n104, S => A(18), Z => n69);
   U101 : NAND3_X1 port map( A1 => n70, A2 => n15, A3 => n69, ZN => p(18));
   U102 : MUX2_X1 port map( A => n100, B => n23, S => A(18), Z => n72);
   U103 : MUX2_X1 port map( A => n99, B => n104, S => A(19), Z => n71);
   U104 : NAND3_X1 port map( A1 => n72, A2 => n15, A3 => n71, ZN => p(19));
   U105 : MUX2_X1 port map( A => n100, B => n101, S => A(19), Z => n74);
   U106 : MUX2_X1 port map( A => n99, B => n95, S => A(20), Z => n73);
   U107 : NAND3_X1 port map( A1 => n74, A2 => n15, A3 => n73, ZN => p(20));
   U108 : MUX2_X1 port map( A => n100, B => n101, S => A(20), Z => n76);
   U109 : MUX2_X1 port map( A => n99, B => n95, S => A(21), Z => n75);
   U110 : NAND3_X1 port map( A1 => n76, A2 => n15, A3 => n75, ZN => p(21));
   U111 : MUX2_X1 port map( A => n100, B => n23, S => A(21), Z => n78);
   U112 : MUX2_X1 port map( A => n99, B => n104, S => A(22), Z => n77);
   U113 : NAND3_X1 port map( A1 => n78, A2 => n15, A3 => n77, ZN => p(22));
   U114 : MUX2_X1 port map( A => n100, B => n23, S => A(22), Z => n80);
   U115 : MUX2_X1 port map( A => n99, B => n95, S => A(23), Z => n79);
   U116 : NAND3_X1 port map( A1 => n80, A2 => n15, A3 => n79, ZN => p(23));
   U117 : MUX2_X1 port map( A => n100, B => n23, S => A(23), Z => n82);
   U118 : MUX2_X1 port map( A => n99, B => n104, S => n105, Z => n81);
   U119 : NAND3_X1 port map( A1 => n82, A2 => n15, A3 => n81, ZN => p(24));
   U120 : MUX2_X1 port map( A => n100, B => n23, S => n105, Z => n84);
   U121 : MUX2_X1 port map( A => n99, B => n104, S => n105, Z => n83);
   U122 : NAND3_X1 port map( A1 => n84, A2 => n97, A3 => n83, ZN => p(25));
   U39 : INV_X1 port map( A => b(0), ZN => n32);
   U10 : BUF_X1 port map( A => n4, Z => n23);
   U4 : CLKBUF_X1 port map( A => n97, Z => n16);
   U13 : BUF_X1 port map( A => n95, Z => n104);
   U14 : INV_X1 port map( A => b(1), ZN => n31);
   n105 <= '0';
   U5 : NAND3_X2 port map( A1 => b(2), A2 => n32, A3 => n31, ZN => n100);
   U6 : CLKBUF_X3 port map( A => n97, Z => n15);
   U7 : OR2_X2 port map( A1 => b(2), A2 => n27, ZN => n95);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_7 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_7;

architecture SYN_beh of ENC_7 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73
      , n74, n75, n76, n77, n78, n79, n86, n88, n90, n91, n92, n93, n94 : 
      std_logic;

begin
   
   U22 : XNOR2_X1 port map( A => b(1), B => b(0), ZN => n17);
   U25 : INV_X1 port map( A => b(2), ZN => n21);
   U27 : INV_X1 port map( A => b(0), ZN => n20);
   U28 : INV_X1 port map( A => b(1), ZN => n19);
   U30 : NAND2_X1 port map( A1 => b(2), A2 => n25, ZN => n22);
   U31 : MUX2_X1 port map( A => n22, B => n86, S => A(0), Z => n18);
   U32 : OAI211_X1 port map( C1 => n21, C2 => n25, A => n91, B => n18, ZN => 
                           p(0));
   U33 : MUX2_X1 port map( A => n91, B => n25, S => A(0), Z => n24);
   U34 : NAND2_X1 port map( A1 => n20, A2 => n19, ZN => n46);
   U36 : NAND4_X1 port map( A1 => n22, A2 => n46, A3 => n92, A4 => n86, ZN => 
                           n88);
   U38 : MUX2_X1 port map( A => n90, B => n86, S => A(1), Z => n23);
   U39 : NAND3_X1 port map( A1 => n24, A2 => n7, A3 => n23, ZN => p(1));
   U40 : MUX2_X1 port map( A => n90, B => n86, S => A(2), Z => n27);
   U41 : MUX2_X1 port map( A => n91, B => n25, S => A(1), Z => n26);
   U42 : NAND3_X1 port map( A1 => n27, A2 => n93, A3 => n26, ZN => p(2));
   U43 : MUX2_X1 port map( A => n91, B => n92, S => A(2), Z => n29);
   U44 : MUX2_X1 port map( A => n90, B => n86, S => A(3), Z => n28);
   U45 : NAND3_X1 port map( A1 => n29, A2 => n93, A3 => n28, ZN => p(3));
   U46 : MUX2_X1 port map( A => n91, B => n92, S => A(3), Z => n31);
   U47 : MUX2_X1 port map( A => n90, B => n86, S => A(4), Z => n30);
   U48 : NAND3_X1 port map( A1 => n31, A2 => n7, A3 => n30, ZN => p(4));
   U49 : MUX2_X1 port map( A => n90, B => n86, S => A(5), Z => n33);
   U50 : MUX2_X1 port map( A => n91, B => n92, S => A(4), Z => n32);
   U51 : NAND3_X1 port map( A1 => n33, A2 => n7, A3 => n32, ZN => p(5));
   U52 : MUX2_X1 port map( A => n91, B => n92, S => A(5), Z => n35);
   U53 : MUX2_X1 port map( A => n90, B => n86, S => A(6), Z => n34);
   U54 : NAND3_X1 port map( A1 => n35, A2 => n93, A3 => n34, ZN => p(6));
   U55 : MUX2_X1 port map( A => n91, B => n92, S => A(6), Z => n37);
   U56 : MUX2_X1 port map( A => n90, B => n86, S => A(7), Z => n36);
   U57 : NAND3_X1 port map( A1 => n37, A2 => n93, A3 => n36, ZN => p(7));
   U58 : MUX2_X1 port map( A => n90, B => n86, S => A(8), Z => n39);
   U59 : MUX2_X1 port map( A => n91, B => n92, S => A(7), Z => n38);
   U60 : NAND3_X1 port map( A1 => n39, A2 => n93, A3 => n38, ZN => p(8));
   U61 : MUX2_X1 port map( A => n91, B => n92, S => A(8), Z => n41);
   U62 : MUX2_X1 port map( A => n90, B => n86, S => A(9), Z => n40);
   U63 : NAND3_X1 port map( A1 => n41, A2 => n7, A3 => n40, ZN => p(9));
   U64 : MUX2_X1 port map( A => n90, B => n86, S => A(10), Z => n43);
   U65 : MUX2_X1 port map( A => n91, B => n92, S => A(9), Z => n42);
   U66 : NAND3_X1 port map( A1 => n93, A2 => n43, A3 => n42, ZN => p(10));
   U67 : MUX2_X1 port map( A => n91, B => n92, S => A(10), Z => n45);
   U68 : MUX2_X1 port map( A => n90, B => n86, S => A(11), Z => n44);
   U69 : NAND3_X1 port map( A1 => n45, A2 => n93, A3 => n44, ZN => p(11));
   U70 : MUX2_X1 port map( A => n91, B => n92, S => A(11), Z => n49);
   U71 : NAND2_X1 port map( A1 => b(2), A2 => n46, ZN => n47);
   U72 : MUX2_X1 port map( A => n47, B => n86, S => A(12), Z => n48);
   U73 : NAND3_X1 port map( A1 => n49, A2 => n7, A3 => n48, ZN => p(12));
   U74 : MUX2_X1 port map( A => n91, B => n92, S => A(12), Z => n51);
   U75 : MUX2_X1 port map( A => n90, B => n86, S => A(13), Z => n50);
   U76 : NAND3_X1 port map( A1 => n51, A2 => n93, A3 => n50, ZN => p(13));
   U77 : MUX2_X1 port map( A => n91, B => n92, S => A(13), Z => n53);
   U78 : MUX2_X1 port map( A => n90, B => n86, S => A(14), Z => n52);
   U79 : NAND3_X1 port map( A1 => n53, A2 => n7, A3 => n52, ZN => p(14));
   U80 : MUX2_X1 port map( A => n91, B => n92, S => A(14), Z => n55);
   U81 : MUX2_X1 port map( A => n90, B => n86, S => A(15), Z => n54);
   U82 : NAND3_X1 port map( A1 => n55, A2 => n93, A3 => n54, ZN => p(15));
   U83 : MUX2_X1 port map( A => n91, B => n92, S => A(15), Z => n57);
   U84 : MUX2_X1 port map( A => n90, B => n86, S => A(16), Z => n56);
   U85 : NAND3_X1 port map( A1 => n57, A2 => n93, A3 => n56, ZN => p(16));
   U86 : MUX2_X1 port map( A => n91, B => n92, S => A(16), Z => n59);
   U87 : MUX2_X1 port map( A => n90, B => n86, S => A(17), Z => n58);
   U88 : NAND3_X1 port map( A1 => n59, A2 => n93, A3 => n58, ZN => p(17));
   U89 : MUX2_X1 port map( A => n91, B => n92, S => A(17), Z => n61);
   U90 : MUX2_X1 port map( A => n90, B => n86, S => A(18), Z => n60);
   U91 : NAND3_X1 port map( A1 => n61, A2 => n93, A3 => n60, ZN => p(18));
   U92 : MUX2_X1 port map( A => n91, B => n92, S => A(18), Z => n63);
   U93 : MUX2_X1 port map( A => n90, B => n86, S => A(19), Z => n62);
   U94 : NAND3_X1 port map( A1 => n63, A2 => n93, A3 => n62, ZN => p(19));
   U95 : MUX2_X1 port map( A => n91, B => n92, S => A(19), Z => n65);
   U96 : MUX2_X1 port map( A => n90, B => n86, S => A(20), Z => n64);
   U97 : NAND3_X1 port map( A1 => n65, A2 => n7, A3 => n64, ZN => p(20));
   U98 : MUX2_X1 port map( A => n91, B => n92, S => A(20), Z => n67);
   U99 : MUX2_X1 port map( A => n90, B => n86, S => A(21), Z => n66);
   U100 : NAND3_X1 port map( A1 => n67, A2 => n7, A3 => n66, ZN => p(21));
   U101 : MUX2_X1 port map( A => n91, B => n92, S => A(21), Z => n69);
   U102 : MUX2_X1 port map( A => n90, B => n86, S => A(22), Z => n68);
   U103 : NAND3_X1 port map( A1 => n69, A2 => n7, A3 => n68, ZN => p(22));
   U104 : MUX2_X1 port map( A => n91, B => n92, S => A(22), Z => n71);
   U105 : MUX2_X1 port map( A => n90, B => n86, S => A(23), Z => n70);
   U106 : NAND3_X1 port map( A1 => n71, A2 => n7, A3 => n70, ZN => p(23));
   U107 : MUX2_X1 port map( A => n91, B => n92, S => A(23), Z => n73);
   U108 : MUX2_X1 port map( A => n90, B => n86, S => n94, Z => n72);
   U109 : NAND3_X1 port map( A1 => n73, A2 => n7, A3 => n72, ZN => p(24));
   U110 : MUX2_X1 port map( A => n91, B => n92, S => n94, Z => n75);
   U111 : MUX2_X1 port map( A => n90, B => n86, S => n94, Z => n74);
   U112 : NAND3_X1 port map( A1 => n75, A2 => n7, A3 => n74, ZN => p(25));
   U113 : MUX2_X1 port map( A => n91, B => n92, S => n94, Z => n77);
   U114 : MUX2_X1 port map( A => n90, B => n86, S => n94, Z => n76);
   U115 : NAND3_X1 port map( A1 => n77, A2 => n7, A3 => n76, ZN => p(26));
   U116 : MUX2_X1 port map( A => n91, B => n92, S => n94, Z => n79);
   U117 : MUX2_X1 port map( A => n90, B => n86, S => n94, Z => n78);
   U118 : NAND3_X1 port map( A1 => n79, A2 => n7, A3 => n78, ZN => p(27));
   U26 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n25);
   U3 : OR2_X2 port map( A1 => b(2), A2 => n17, ZN => n86);
   U29 : NAND3_X1 port map( A1 => b(2), A2 => n20, A3 => n19, ZN => n91);
   U4 : BUF_X2 port map( A => n88, Z => n7);
   U5 : BUF_X1 port map( A => n88, Z => n93);
   n94 <= '0';
   U6 : NAND3_X2 port map( A1 => b(1), A2 => n21, A3 => b(0), ZN => n92);
   U8 : NAND2_X2 port map( A1 => b(2), A2 => n46, ZN => n90);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_8 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_8;

architecture SYN_beh of ENC_8 is

   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
      n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44
      , n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, 
      n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73
      , n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n86, n88, n90, n91, 
      n92, n96 : std_logic;

begin
   
   U18 : XNOR2_X1 port map( A => b(1), B => b(0), ZN => n16);
   U22 : INV_X1 port map( A => b(2), ZN => n19);
   U23 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n18);
   U24 : INV_X1 port map( A => b(0), ZN => n22);
   U25 : INV_X1 port map( A => b(1), ZN => n21);
   U27 : NAND2_X1 port map( A1 => b(2), A2 => n18, ZN => n20);
   U28 : MUX2_X1 port map( A => n20, B => n86, S => A(0), Z => n17);
   U29 : OAI211_X1 port map( C1 => n19, C2 => n18, A => n91, B => n17, ZN => 
                           p(0));
   U31 : MUX2_X1 port map( A => n91, B => n92, S => A(0), Z => n24);
   U33 : NAND2_X1 port map( A1 => n22, A2 => n21, ZN => n45);
   U35 : MUX2_X1 port map( A => n90, B => n86, S => A(1), Z => n23);
   U36 : NAND3_X1 port map( A1 => n24, A2 => n88, A3 => n23, ZN => p(1));
   U37 : MUX2_X1 port map( A => n91, B => n92, S => A(1), Z => n26);
   U38 : MUX2_X1 port map( A => n90, B => n86, S => A(2), Z => n25);
   U39 : NAND3_X1 port map( A1 => n26, A2 => n88, A3 => n25, ZN => p(2));
   U40 : MUX2_X1 port map( A => n91, B => n92, S => A(2), Z => n28);
   U41 : MUX2_X1 port map( A => n90, B => n86, S => A(3), Z => n27);
   U42 : NAND3_X1 port map( A1 => n28, A2 => n88, A3 => n27, ZN => p(3));
   U43 : MUX2_X1 port map( A => n91, B => n92, S => A(3), Z => n30);
   U44 : MUX2_X1 port map( A => n90, B => n86, S => A(4), Z => n29);
   U45 : NAND3_X1 port map( A1 => n30, A2 => n88, A3 => n29, ZN => p(4));
   U46 : MUX2_X1 port map( A => n91, B => n92, S => A(4), Z => n32);
   U47 : MUX2_X1 port map( A => n90, B => n86, S => A(5), Z => n31);
   U48 : NAND3_X1 port map( A1 => n31, A2 => n88, A3 => n32, ZN => p(5));
   U49 : MUX2_X1 port map( A => n91, B => n92, S => A(5), Z => n34);
   U50 : MUX2_X1 port map( A => n90, B => n86, S => A(6), Z => n33);
   U51 : NAND3_X1 port map( A1 => n34, A2 => n88, A3 => n33, ZN => p(6));
   U52 : NAND2_X1 port map( A1 => b(2), A2 => n45, ZN => n52);
   U53 : MUX2_X1 port map( A => n52, B => n86, S => A(7), Z => n36);
   U54 : MUX2_X1 port map( A => n91, B => n92, S => A(6), Z => n35);
   U55 : NAND3_X1 port map( A1 => n36, A2 => n88, A3 => n35, ZN => p(7));
   U56 : MUX2_X1 port map( A => n90, B => n86, S => A(8), Z => n38);
   U57 : MUX2_X1 port map( A => n91, B => n92, S => A(7), Z => n37);
   U58 : NAND3_X1 port map( A1 => n38, A2 => n88, A3 => n37, ZN => p(8));
   U59 : MUX2_X1 port map( A => n91, B => n92, S => A(8), Z => n40);
   U60 : MUX2_X1 port map( A => n90, B => n86, S => A(9), Z => n39);
   U61 : NAND3_X1 port map( A1 => n40, A2 => n88, A3 => n39, ZN => p(9));
   U62 : MUX2_X1 port map( A => n91, B => n92, S => A(9), Z => n42);
   U63 : MUX2_X1 port map( A => n90, B => n86, S => A(10), Z => n41);
   U64 : NAND3_X1 port map( A1 => n42, A2 => n88, A3 => n41, ZN => p(10));
   U65 : MUX2_X1 port map( A => n91, B => n92, S => A(10), Z => n44);
   U66 : MUX2_X1 port map( A => n90, B => n86, S => A(11), Z => n43);
   U67 : NAND3_X1 port map( A1 => n44, A2 => n88, A3 => n43, ZN => p(11));
   U68 : MUX2_X1 port map( A => n91, B => n92, S => A(11), Z => n47);
   U69 : NAND2_X1 port map( A1 => b(2), A2 => n45, ZN => n63);
   U70 : MUX2_X1 port map( A => n63, B => n86, S => A(12), Z => n46);
   U71 : NAND3_X1 port map( A1 => n47, A2 => n88, A3 => n46, ZN => p(12));
   U72 : MUX2_X1 port map( A => n52, B => n86, S => A(13), Z => n49);
   U73 : MUX2_X1 port map( A => n91, B => n92, S => A(12), Z => n48);
   U74 : NAND3_X1 port map( A1 => n49, A2 => n48, A3 => n88, ZN => p(13));
   U75 : MUX2_X1 port map( A => n91, B => n92, S => A(13), Z => n51);
   U76 : MUX2_X1 port map( A => n52, B => n86, S => A(14), Z => n50);
   U77 : NAND3_X1 port map( A1 => n51, A2 => n88, A3 => n50, ZN => p(14));
   U78 : MUX2_X1 port map( A => n52, B => n86, S => A(15), Z => n54);
   U79 : MUX2_X1 port map( A => n91, B => n92, S => A(14), Z => n53);
   U80 : NAND3_X1 port map( A1 => n54, A2 => n53, A3 => n88, ZN => p(15));
   U81 : MUX2_X1 port map( A => n91, B => n92, S => A(15), Z => n56);
   U82 : MUX2_X1 port map( A => n63, B => n86, S => A(16), Z => n55);
   U83 : NAND3_X1 port map( A1 => n56, A2 => n88, A3 => n55, ZN => p(16));
   U84 : MUX2_X1 port map( A => n63, B => n86, S => A(17), Z => n58);
   U85 : MUX2_X1 port map( A => n91, B => n92, S => A(16), Z => n57);
   U86 : NAND3_X1 port map( A1 => n58, A2 => n57, A3 => n88, ZN => p(17));
   U87 : MUX2_X1 port map( A => n91, B => n92, S => A(17), Z => n60);
   U88 : MUX2_X1 port map( A => n90, B => n86, S => A(18), Z => n59);
   U89 : NAND3_X1 port map( A1 => n60, A2 => n88, A3 => n59, ZN => p(18));
   U90 : MUX2_X1 port map( A => n63, B => n86, S => A(19), Z => n62);
   U91 : MUX2_X1 port map( A => n91, B => n92, S => A(18), Z => n61);
   U92 : NAND3_X1 port map( A1 => n62, A2 => n61, A3 => n88, ZN => p(19));
   U93 : MUX2_X1 port map( A => n63, B => n86, S => A(20), Z => n65);
   U94 : MUX2_X1 port map( A => n91, B => n92, S => A(19), Z => n64);
   U95 : NAND3_X1 port map( A1 => n88, A2 => n65, A3 => n64, ZN => p(20));
   U96 : MUX2_X1 port map( A => n91, B => n92, S => A(20), Z => n67);
   U97 : MUX2_X1 port map( A => n90, B => n86, S => A(21), Z => n66);
   U98 : NAND3_X1 port map( A1 => n67, A2 => n88, A3 => n66, ZN => p(21));
   U99 : MUX2_X1 port map( A => n91, B => n92, S => A(21), Z => n69);
   U100 : MUX2_X1 port map( A => n90, B => n86, S => A(22), Z => n68);
   U101 : NAND3_X1 port map( A1 => n69, A2 => n88, A3 => n68, ZN => p(22));
   U102 : MUX2_X1 port map( A => n91, B => n92, S => A(22), Z => n71);
   U103 : MUX2_X1 port map( A => n90, B => n86, S => A(23), Z => n70);
   U104 : NAND3_X1 port map( A1 => n71, A2 => n88, A3 => n70, ZN => p(23));
   U105 : MUX2_X1 port map( A => n91, B => n92, S => A(23), Z => n73);
   U106 : MUX2_X1 port map( A => n90, B => n86, S => n96, Z => n72);
   U107 : NAND3_X1 port map( A1 => n73, A2 => n88, A3 => n72, ZN => p(24));
   U108 : MUX2_X1 port map( A => n91, B => n92, S => n96, Z => n75);
   U109 : MUX2_X1 port map( A => n90, B => n86, S => n96, Z => n74);
   U110 : NAND3_X1 port map( A1 => n75, A2 => n88, A3 => n74, ZN => p(25));
   U111 : MUX2_X1 port map( A => n91, B => n92, S => n96, Z => n77);
   U112 : MUX2_X1 port map( A => n90, B => n86, S => n96, Z => n76);
   U113 : NAND3_X1 port map( A1 => n77, A2 => n88, A3 => n76, ZN => p(26));
   U114 : MUX2_X1 port map( A => n91, B => n92, S => n96, Z => n79);
   U115 : MUX2_X1 port map( A => n90, B => n86, S => n96, Z => n78);
   U116 : NAND3_X1 port map( A1 => n79, A2 => n88, A3 => n78, ZN => p(27));
   U117 : MUX2_X1 port map( A => n91, B => n92, S => n96, Z => n81);
   U118 : MUX2_X1 port map( A => n90, B => n86, S => n96, Z => n80);
   U119 : NAND3_X1 port map( A1 => n81, A2 => n88, A3 => n80, ZN => p(28));
   U120 : MUX2_X1 port map( A => n91, B => n92, S => n96, Z => n83);
   U121 : MUX2_X1 port map( A => n90, B => n86, S => n96, Z => n82);
   U122 : NAND3_X1 port map( A1 => n83, A2 => n88, A3 => n82, ZN => p(29));
   U32 : NAND2_X2 port map( A1 => b(2), A2 => n20, ZN => n88);
   U26 : NAND3_X1 port map( A1 => b(2), A2 => n22, A3 => n21, ZN => n91);
   U34 : NAND2_X1 port map( A1 => b(2), A2 => n45, ZN => n90);
   U4 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n92);
   n96 <= '0';
   U3 : OR2_X2 port map( A1 => b(2), A2 => n16, ZN => n86);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_9 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_9;

architecture SYN_beh of ENC_9 is

   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
      n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n104 : std_logic;

begin
   
   U5 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n32);
   U14 : NAND4_X1 port map( A1 => n31, A2 => n32, A3 => n99, A4 => n93, ZN => 
                           n6);
   U26 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n25);
   U30 : INV_X1 port map( A => b(2), ZN => n28);
   U31 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n27);
   U32 : INV_X1 port map( A => b(0), ZN => n30);
   U33 : INV_X1 port map( A => b(1), ZN => n29);
   U35 : NAND2_X1 port map( A1 => b(2), A2 => n27, ZN => n31);
   U36 : MUX2_X1 port map( A => n31, B => n93, S => A(0), Z => n26);
   U37 : OAI211_X1 port map( C1 => n28, C2 => n27, A => n98, B => n26, ZN => 
                           p(0));
   U39 : MUX2_X1 port map( A => n98, B => n99, S => A(0), Z => n34);
   U40 : NAND4_X1 port map( A1 => n31, A2 => n32, A3 => n99, A4 => n93, ZN => 
                           n95);
   U42 : MUX2_X1 port map( A => n97, B => n93, S => A(1), Z => n33);
   U43 : NAND3_X1 port map( A1 => n34, A2 => n95, A3 => n33, ZN => p(1));
   U44 : MUX2_X1 port map( A => n98, B => n99, S => A(1), Z => n36);
   U45 : MUX2_X1 port map( A => n97, B => n93, S => A(2), Z => n35);
   U46 : NAND3_X1 port map( A1 => n36, A2 => n95, A3 => n35, ZN => p(2));
   U47 : MUX2_X1 port map( A => n98, B => n99, S => A(2), Z => n38);
   U48 : MUX2_X1 port map( A => n97, B => n93, S => A(3), Z => n37);
   U49 : NAND3_X1 port map( A1 => n38, A2 => n95, A3 => n37, ZN => p(3));
   U50 : MUX2_X1 port map( A => n98, B => n99, S => A(3), Z => n40);
   U51 : MUX2_X1 port map( A => n97, B => n93, S => A(4), Z => n39);
   U52 : NAND3_X1 port map( A1 => n40, A2 => n5, A3 => n39, ZN => p(4));
   U53 : MUX2_X1 port map( A => n98, B => n99, S => A(4), Z => n42);
   U54 : MUX2_X1 port map( A => n97, B => n93, S => A(5), Z => n41);
   U55 : NAND3_X1 port map( A1 => n42, A2 => n5, A3 => n41, ZN => p(5));
   U56 : MUX2_X1 port map( A => n98, B => n99, S => A(5), Z => n44);
   U57 : MUX2_X1 port map( A => n97, B => n93, S => A(6), Z => n43);
   U58 : NAND3_X1 port map( A1 => n44, A2 => n95, A3 => n43, ZN => p(6));
   U59 : MUX2_X1 port map( A => n98, B => n99, S => A(6), Z => n46);
   U60 : MUX2_X1 port map( A => n97, B => n93, S => A(7), Z => n45);
   U61 : NAND3_X1 port map( A1 => n46, A2 => n95, A3 => n45, ZN => p(7));
   U62 : MUX2_X1 port map( A => n98, B => n99, S => A(7), Z => n48);
   U63 : MUX2_X1 port map( A => n97, B => n93, S => A(8), Z => n47);
   U64 : NAND3_X1 port map( A1 => n47, A2 => n6, A3 => n48, ZN => p(8));
   U65 : MUX2_X1 port map( A => n98, B => n99, S => A(8), Z => n50);
   U66 : MUX2_X1 port map( A => n97, B => n93, S => A(9), Z => n49);
   U67 : NAND3_X1 port map( A1 => n50, A2 => n5, A3 => n49, ZN => p(9));
   U68 : MUX2_X1 port map( A => n98, B => n99, S => A(9), Z => n52);
   U69 : MUX2_X1 port map( A => n97, B => n93, S => A(10), Z => n51);
   U70 : NAND3_X1 port map( A1 => n52, A2 => n95, A3 => n51, ZN => p(10));
   U71 : MUX2_X1 port map( A => n97, B => n93, S => A(11), Z => n54);
   U72 : MUX2_X1 port map( A => n98, B => n99, S => A(10), Z => n53);
   U73 : NAND3_X1 port map( A1 => n54, A2 => n5, A3 => n53, ZN => p(11));
   U74 : MUX2_X1 port map( A => n98, B => n99, S => A(11), Z => n56);
   U75 : MUX2_X1 port map( A => n97, B => n93, S => A(12), Z => n55);
   U76 : NAND3_X1 port map( A1 => n56, A2 => n5, A3 => n55, ZN => p(12));
   U77 : MUX2_X1 port map( A => n98, B => n99, S => A(12), Z => n58);
   U78 : MUX2_X1 port map( A => n97, B => n93, S => A(13), Z => n57);
   U79 : NAND3_X1 port map( A1 => n58, A2 => n6, A3 => n57, ZN => p(13));
   U80 : MUX2_X1 port map( A => n98, B => n99, S => A(13), Z => n60);
   U81 : MUX2_X1 port map( A => n97, B => n93, S => A(14), Z => n59);
   U82 : NAND3_X1 port map( A1 => n60, A2 => n5, A3 => n59, ZN => p(14));
   U83 : MUX2_X1 port map( A => n98, B => n99, S => A(14), Z => n62);
   U84 : MUX2_X1 port map( A => n97, B => n93, S => A(15), Z => n61);
   U85 : NAND3_X1 port map( A1 => n62, A2 => n95, A3 => n61, ZN => p(15));
   U86 : MUX2_X1 port map( A => n98, B => n99, S => A(15), Z => n64);
   U87 : MUX2_X1 port map( A => n97, B => n93, S => A(16), Z => n63);
   U88 : NAND3_X1 port map( A1 => n64, A2 => n5, A3 => n63, ZN => p(16));
   U89 : MUX2_X1 port map( A => n97, B => n93, S => A(17), Z => n66);
   U90 : MUX2_X1 port map( A => n98, B => n99, S => A(16), Z => n65);
   U91 : NAND3_X1 port map( A1 => n66, A2 => n5, A3 => n65, ZN => p(17));
   U92 : MUX2_X1 port map( A => n98, B => n99, S => A(17), Z => n68);
   U93 : MUX2_X1 port map( A => n97, B => n93, S => A(18), Z => n67);
   U94 : NAND3_X1 port map( A1 => n68, A2 => n5, A3 => n67, ZN => p(18));
   U95 : MUX2_X1 port map( A => n98, B => n99, S => A(18), Z => n70);
   U96 : MUX2_X1 port map( A => n97, B => n93, S => A(19), Z => n69);
   U97 : NAND3_X1 port map( A1 => n70, A2 => n95, A3 => n69, ZN => p(19));
   U98 : MUX2_X1 port map( A => n98, B => n99, S => A(19), Z => n72);
   U99 : MUX2_X1 port map( A => n97, B => n93, S => A(20), Z => n71);
   U100 : NAND3_X1 port map( A1 => n72, A2 => n6, A3 => n71, ZN => p(20));
   U101 : MUX2_X1 port map( A => n97, B => n93, S => A(21), Z => n74);
   U102 : MUX2_X1 port map( A => n98, B => n99, S => A(20), Z => n73);
   U103 : NAND3_X1 port map( A1 => n74, A2 => n5, A3 => n73, ZN => p(21));
   U104 : MUX2_X1 port map( A => n97, B => n93, S => A(22), Z => n76);
   U105 : MUX2_X1 port map( A => n98, B => n99, S => A(21), Z => n75);
   U106 : NAND3_X1 port map( A1 => n6, A2 => n76, A3 => n75, ZN => p(22));
   U107 : MUX2_X1 port map( A => n98, B => n99, S => A(22), Z => n78);
   U108 : MUX2_X1 port map( A => n97, B => n93, S => A(23), Z => n77);
   U109 : NAND3_X1 port map( A1 => n78, A2 => n5, A3 => n77, ZN => p(23));
   U110 : MUX2_X1 port map( A => n98, B => n99, S => A(23), Z => n80);
   U111 : MUX2_X1 port map( A => n97, B => n93, S => n104, Z => n79);
   U112 : NAND3_X1 port map( A1 => n80, A2 => n5, A3 => n79, ZN => p(24));
   U113 : MUX2_X1 port map( A => n98, B => n99, S => n104, Z => n82);
   U114 : MUX2_X1 port map( A => n97, B => n93, S => n104, Z => n81);
   U115 : NAND3_X1 port map( A1 => n82, A2 => n6, A3 => n81, ZN => p(25));
   U116 : MUX2_X1 port map( A => n98, B => n99, S => n104, Z => n84);
   U117 : MUX2_X1 port map( A => n97, B => n93, S => n104, Z => n83);
   U118 : NAND3_X1 port map( A1 => n84, A2 => n5, A3 => n83, ZN => p(26));
   U119 : MUX2_X1 port map( A => n98, B => n99, S => n104, Z => n86);
   U120 : MUX2_X1 port map( A => n97, B => n93, S => n104, Z => n85);
   U121 : NAND3_X1 port map( A1 => n86, A2 => n95, A3 => n85, ZN => p(27));
   U122 : MUX2_X1 port map( A => n98, B => n99, S => n104, Z => n88);
   U123 : MUX2_X1 port map( A => n97, B => n93, S => n104, Z => n87);
   U124 : NAND3_X1 port map( A1 => n88, A2 => n5, A3 => n87, ZN => p(28));
   U125 : MUX2_X1 port map( A => n98, B => n99, S => n104, Z => n90);
   U126 : MUX2_X1 port map( A => n97, B => n93, S => n104, Z => n89);
   U127 : NAND3_X1 port map( A1 => n90, A2 => n95, A3 => n89, ZN => p(29));
   U128 : MUX2_X1 port map( A => n98, B => n99, S => n104, Z => n92);
   U129 : MUX2_X1 port map( A => n97, B => n93, S => n104, Z => n91);
   U130 : NAND3_X1 port map( A1 => n92, A2 => n6, A3 => n91, ZN => p(30));
   U131 : MUX2_X1 port map( A => n98, B => n99, S => n104, Z => n96);
   U132 : MUX2_X1 port map( A => n97, B => n93, S => n104, Z => n94);
   U133 : NAND3_X1 port map( A1 => n96, A2 => n95, A3 => n94, ZN => p(31));
   U13 : NAND4_X1 port map( A1 => n32, A2 => n93, A3 => n31, A4 => n99, ZN => 
                           n5);
   U34 : NAND3_X1 port map( A1 => b(2), A2 => n30, A3 => n29, ZN => n98);
   U41 : NAND2_X2 port map( A1 => b(2), A2 => n32, ZN => n97);
   U6 : OR2_X2 port map( A1 => n25, A2 => b(2), ZN => n93);
   n104 <= '0';
   U3 : NAND3_X2 port map( A1 => b(0), A2 => n28, A3 => b(1), ZN => n99);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_10 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_10;

architecture SYN_beh of ENC_10 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n9, n10, n11, n12, n13, n14, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n108, n110, n111 : std_logic;

begin
   
   U5 : AND3_X1 port map( A1 => b(2), A2 => n30, A3 => n29, ZN => n12);
   U6 : XNOR2_X1 port map( A => b(0), B => n29, ZN => n10);
   U10 : NAND2_X1 port map( A1 => n30, A2 => n29, ZN => n69);
   U13 : NAND2_X1 port map( A1 => n80, A2 => n3, ZN => n4);
   U14 : NAND2_X1 port map( A1 => n89, A2 => A(16), ZN => n5);
   U15 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => n64);
   U16 : INV_X1 port map( A => A(16), ZN => n3);
   U22 : NAND2_X1 port map( A1 => n10, A2 => n58, ZN => n102);
   U26 : NAND2_X1 port map( A1 => n69, A2 => n58, ZN => n13);
   U27 : NAND2_X1 port map( A1 => n10, A2 => n58, ZN => n14);
   U32 : INV_X1 port map( A => A(18), ZN => n27);
   U33 : INV_X1 port map( A => b(2), ZN => n58);
   U37 : NAND2_X1 port map( A1 => b(2), A2 => n65, ZN => n31);
   U38 : MUX2_X1 port map( A => n31, B => n14, S => A(0), Z => n28);
   U39 : OAI211_X1 port map( C1 => n58, C2 => n65, A => n28, B => n110, ZN => 
                           p(0));
   U40 : MUX2_X1 port map( A => n110, B => n65, S => A(0), Z => n33);
   U41 : NAND2_X1 port map( A1 => n69, A2 => n58, ZN => n72);
   U43 : MUX2_X1 port map( A => n106, B => n102, S => A(1), Z => n32);
   U44 : NAND3_X1 port map( A1 => n33, A2 => n108, A3 => n32, ZN => p(1));
   U45 : MUX2_X1 port map( A => n110, B => n65, S => A(1), Z => n35);
   U46 : MUX2_X1 port map( A => n106, B => n14, S => A(2), Z => n34);
   U47 : NAND3_X1 port map( A1 => n35, A2 => n108, A3 => n34, ZN => p(2));
   U48 : MUX2_X1 port map( A => n110, B => n65, S => A(2), Z => n37);
   U49 : MUX2_X1 port map( A => n106, B => n102, S => A(3), Z => n36);
   U50 : NAND3_X1 port map( A1 => n37, A2 => n108, A3 => n36, ZN => p(3));
   U51 : MUX2_X1 port map( A => n110, B => n65, S => A(3), Z => n39);
   U52 : MUX2_X1 port map( A => n106, B => n14, S => A(4), Z => n38);
   U53 : NAND3_X1 port map( A1 => n39, A2 => n108, A3 => n38, ZN => p(4));
   U54 : MUX2_X1 port map( A => n110, B => n65, S => A(4), Z => n41);
   U55 : MUX2_X1 port map( A => n106, B => n102, S => A(5), Z => n40);
   U56 : NAND3_X1 port map( A1 => n41, A2 => n108, A3 => n40, ZN => p(5));
   U57 : MUX2_X1 port map( A => n110, B => n65, S => A(5), Z => n43);
   U58 : MUX2_X1 port map( A => n106, B => n14, S => A(6), Z => n42);
   U59 : NAND3_X1 port map( A1 => n43, A2 => n108, A3 => n42, ZN => p(6));
   U60 : MUX2_X1 port map( A => n110, B => n65, S => A(6), Z => n45);
   U61 : MUX2_X1 port map( A => n106, B => n102, S => A(7), Z => n44);
   U62 : NAND3_X1 port map( A1 => n45, A2 => n108, A3 => n44, ZN => p(7));
   U63 : MUX2_X1 port map( A => n110, B => n65, S => A(7), Z => n47);
   U64 : MUX2_X1 port map( A => n106, B => n14, S => A(8), Z => n46);
   U65 : NAND3_X1 port map( A1 => n47, A2 => n108, A3 => n46, ZN => p(8));
   U66 : MUX2_X1 port map( A => n110, B => n65, S => A(8), Z => n49);
   U67 : NAND2_X1 port map( A1 => b(2), A2 => n69, ZN => n80);
   U68 : MUX2_X1 port map( A => n80, B => n102, S => A(9), Z => n48);
   U69 : NAND3_X1 port map( A1 => n49, A2 => n108, A3 => n48, ZN => p(9));
   U70 : MUX2_X1 port map( A => n110, B => n65, S => A(9), Z => n51);
   U71 : MUX2_X1 port map( A => n106, B => n14, S => A(10), Z => n50);
   U72 : NAND3_X1 port map( A1 => n51, A2 => n108, A3 => n50, ZN => p(10));
   U73 : MUX2_X1 port map( A => n110, B => n65, S => A(10), Z => n53);
   U74 : MUX2_X1 port map( A => n80, B => n102, S => A(11), Z => n52);
   U75 : NAND3_X1 port map( A1 => n53, A2 => n108, A3 => n52, ZN => p(11));
   U76 : MUX2_X1 port map( A => n110, B => n65, S => A(11), Z => n55);
   U77 : MUX2_X1 port map( A => n106, B => n14, S => A(12), Z => n54);
   U78 : NAND3_X1 port map( A1 => n55, A2 => n108, A3 => n54, ZN => p(12));
   U79 : MUX2_X1 port map( A => n110, B => n65, S => A(12), Z => n57);
   U80 : MUX2_X1 port map( A => n106, B => n102, S => A(13), Z => n56);
   U81 : NAND3_X1 port map( A1 => n57, A2 => n108, A3 => n56, ZN => p(13));
   U82 : NAND2_X1 port map( A1 => n10, A2 => n58, ZN => n89);
   U83 : MUX2_X1 port map( A => n80, B => n89, S => A(14), Z => n60);
   U84 : MUX2_X1 port map( A => n110, B => n65, S => A(13), Z => n59);
   U85 : NAND3_X1 port map( A1 => n60, A2 => n108, A3 => n59, ZN => p(14));
   U86 : MUX2_X1 port map( A => n110, B => n65, S => A(14), Z => n62);
   U87 : MUX2_X1 port map( A => n106, B => n89, S => A(15), Z => n61);
   U88 : NAND3_X1 port map( A1 => n62, A2 => n108, A3 => n61, ZN => p(15));
   U89 : MUX2_X1 port map( A => n110, B => n65, S => A(15), Z => n63);
   U90 : NAND3_X1 port map( A1 => n64, A2 => n63, A3 => n108, ZN => p(16));
   U91 : MUX2_X1 port map( A => n110, B => n65, S => A(16), Z => n68);
   U93 : OAI21_X1 port map( B1 => b(2), B2 => n11, A => A(17), ZN => n66);
   U94 : OAI211_X1 port map( C1 => A(17), C2 => b(2), A => n66, B => n69, ZN =>
                           n67);
   U95 : NAND3_X1 port map( A1 => n68, A2 => n67, A3 => n108, ZN => p(17));
   U96 : INV_X1 port map( A => n69, ZN => n71);
   U97 : INV_X1 port map( A => n13, ZN => n70);
   U98 : OAI33_X1 port map( A1 => n11, A2 => n13, A3 => n27, B1 => A(18), B2 =>
                           n71, B3 => n70, ZN => n75);
   U99 : MUX2_X1 port map( A => n12, B => n11, S => A(17), Z => n74);
   U100 : OR3_X1 port map( A1 => n9, A2 => n75, A3 => n74, ZN => p(18));
   U101 : MUX2_X1 port map( A => n110, B => n65, S => A(18), Z => n77);
   U102 : MUX2_X1 port map( A => n80, B => n89, S => A(19), Z => n76);
   U103 : NAND3_X1 port map( A1 => n77, A2 => n108, A3 => n76, ZN => p(19));
   U104 : MUX2_X1 port map( A => n110, B => n65, S => A(19), Z => n79);
   U105 : MUX2_X1 port map( A => n80, B => n89, S => A(20), Z => n78);
   U106 : NAND3_X1 port map( A1 => n79, A2 => n108, A3 => n78, ZN => p(20));
   U107 : MUX2_X1 port map( A => n110, B => n65, S => A(20), Z => n82);
   U108 : MUX2_X1 port map( A => n80, B => n89, S => A(21), Z => n81);
   U109 : NAND3_X1 port map( A1 => n82, A2 => n108, A3 => n81, ZN => p(21));
   U110 : MUX2_X1 port map( A => n110, B => n65, S => A(21), Z => n84);
   U111 : MUX2_X1 port map( A => n106, B => n89, S => A(22), Z => n83);
   U112 : NAND3_X1 port map( A1 => n84, A2 => n108, A3 => n83, ZN => p(22));
   U113 : MUX2_X1 port map( A => n110, B => n65, S => A(22), Z => n86);
   U114 : MUX2_X1 port map( A => n106, B => n89, S => A(23), Z => n85);
   U115 : NAND3_X1 port map( A1 => n86, A2 => n108, A3 => n85, ZN => p(23));
   U116 : MUX2_X1 port map( A => n110, B => n65, S => A(23), Z => n88);
   U117 : MUX2_X1 port map( A => n106, B => n102, S => n111, Z => n87);
   U118 : NAND3_X1 port map( A1 => n88, A2 => n108, A3 => n87, ZN => p(24));
   U119 : MUX2_X1 port map( A => n110, B => n65, S => n111, Z => n91);
   U120 : MUX2_X1 port map( A => n106, B => n14, S => n111, Z => n90);
   U121 : NAND3_X1 port map( A1 => n91, A2 => n108, A3 => n90, ZN => p(25));
   U122 : MUX2_X1 port map( A => n110, B => n65, S => n111, Z => n93);
   U123 : MUX2_X1 port map( A => n106, B => n14, S => n111, Z => n92);
   U124 : NAND3_X1 port map( A1 => n93, A2 => n108, A3 => n92, ZN => p(26));
   U125 : MUX2_X1 port map( A => n110, B => n65, S => n111, Z => n95);
   U126 : MUX2_X1 port map( A => n106, B => n102, S => n111, Z => n94);
   U127 : NAND3_X1 port map( A1 => n95, A2 => n108, A3 => n94, ZN => p(27));
   U128 : MUX2_X1 port map( A => n110, B => n65, S => n111, Z => n97);
   U129 : MUX2_X1 port map( A => n106, B => n14, S => n111, Z => n96);
   U130 : NAND3_X1 port map( A1 => n97, A2 => n108, A3 => n96, ZN => p(28));
   U131 : MUX2_X1 port map( A => n110, B => n65, S => n111, Z => n99);
   U132 : MUX2_X1 port map( A => n106, B => n102, S => n111, Z => n98);
   U133 : NAND3_X1 port map( A1 => n99, A2 => n108, A3 => n98, ZN => p(29));
   U134 : MUX2_X1 port map( A => n110, B => n65, S => n111, Z => n101);
   U135 : MUX2_X1 port map( A => n106, B => n14, S => n111, Z => n100);
   U136 : NAND3_X1 port map( A1 => n101, A2 => n108, A3 => n100, ZN => p(30));
   U137 : MUX2_X1 port map( A => n106, B => n102, S => n111, Z => n104);
   U138 : MUX2_X1 port map( A => n110, B => n65, S => n111, Z => n103);
   U139 : NAND3_X1 port map( A1 => n108, A2 => n104, A3 => n103, ZN => p(31));
   U140 : MUX2_X1 port map( A => n110, B => n65, S => n111, Z => n105);
   U141 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => p(32));
   U11 : AND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n11);
   U17 : AND3_X1 port map( A1 => n31, A2 => n69, A3 => n72, ZN => n9);
   U4 : INV_X2 port map( A => n9, ZN => n108);
   U12 : INV_X1 port map( A => b(0), ZN => n30);
   U19 : INV_X1 port map( A => b(1), ZN => n29);
   n111 <= '0';
   U3 : NAND2_X2 port map( A1 => b(1), A2 => b(0), ZN => n65);
   U7 : INV_X2 port map( A => n12, ZN => n110);
   U8 : NAND2_X2 port map( A1 => b(2), A2 => n69, ZN => n106);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_11 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_11;

architecture SYN_beh of ENC_11 is

   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n5, n6, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23
      , n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, 
      n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52
      , n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n93 : std_logic;

begin
   
   U3 : OR2_X1 port map( A1 => n1, A2 => b(2), ZN => n70);
   U4 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n1);
   U7 : NAND2_X1 port map( A1 => b(2), A2 => n24, ZN => n4);
   U8 : NAND2_X1 port map( A1 => b(2), A2 => n24, ZN => n78);
   U15 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => b(2), ZN => n5);
   U17 : NAND3_X1 port map( A1 => b(0), A2 => b(1), A3 => b(2), ZN => n15);
   U19 : INV_X1 port map( A => b(0), ZN => n45);
   U20 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => b(2), ZN => n88);
   U22 : XOR2_X1 port map( A => b(0), B => b(1), Z => n13);
   U23 : NAND2_X1 port map( A1 => n13, A2 => n37, ZN => n83);
   U24 : MUX2_X1 port map( A => n37, B => n6, S => A(0), Z => n14);
   U25 : NAND3_X1 port map( A1 => n15, A2 => n88, A3 => n14, ZN => p(0));
   U27 : MUX2_X1 port map( A => n5, B => n87, S => A(0), Z => n17);
   U29 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => n24);
   U30 : NAND2_X1 port map( A1 => b(2), A2 => n24, ZN => n90);
   U31 : MUX2_X1 port map( A => n4, B => n6, S => A(1), Z => n16);
   U32 : NAND3_X1 port map( A1 => n17, A2 => n85, A3 => n16, ZN => p(1));
   U33 : MUX2_X1 port map( A => n88, B => n87, S => A(1), Z => n19);
   U34 : MUX2_X1 port map( A => n92, B => n6, S => A(2), Z => n18);
   U35 : NAND3_X1 port map( A1 => n19, A2 => n85, A3 => n18, ZN => p(2));
   U36 : MUX2_X1 port map( A => n5, B => n87, S => A(2), Z => n21);
   U37 : MUX2_X1 port map( A => n4, B => n6, S => A(3), Z => n20);
   U38 : NAND3_X1 port map( A1 => n21, A2 => n85, A3 => n20, ZN => p(3));
   U39 : MUX2_X1 port map( A => n88, B => n87, S => A(3), Z => n23);
   U40 : MUX2_X1 port map( A => n4, B => n6, S => A(4), Z => n22);
   U41 : NAND3_X1 port map( A1 => n23, A2 => n85, A3 => n22, ZN => p(4));
   U42 : MUX2_X1 port map( A => n5, B => n87, S => A(4), Z => n26);
   U43 : MUX2_X1 port map( A => n90, B => n6, S => A(5), Z => n25);
   U44 : NAND3_X1 port map( A1 => n26, A2 => n85, A3 => n25, ZN => p(5));
   U45 : MUX2_X1 port map( A => n88, B => n87, S => A(5), Z => n28);
   U46 : MUX2_X1 port map( A => n4, B => n6, S => A(6), Z => n27);
   U47 : NAND3_X1 port map( A1 => n28, A2 => n85, A3 => n27, ZN => p(6));
   U48 : MUX2_X1 port map( A => n5, B => n87, S => A(6), Z => n30);
   U49 : MUX2_X1 port map( A => n92, B => n6, S => A(7), Z => n29);
   U50 : NAND3_X1 port map( A1 => n30, A2 => n85, A3 => n29, ZN => p(7));
   U51 : MUX2_X1 port map( A => n88, B => n87, S => A(7), Z => n32);
   U52 : MUX2_X1 port map( A => n4, B => n83, S => A(8), Z => n31);
   U53 : NAND3_X1 port map( A1 => n32, A2 => n85, A3 => n31, ZN => p(8));
   U54 : MUX2_X1 port map( A => n5, B => n87, S => A(8), Z => n34);
   U55 : MUX2_X1 port map( A => n4, B => n6, S => A(9), Z => n33);
   U56 : NAND3_X1 port map( A1 => n34, A2 => n85, A3 => n33, ZN => p(9));
   U57 : MUX2_X1 port map( A => n90, B => n6, S => A(10), Z => n36);
   U58 : MUX2_X1 port map( A => n88, B => n87, S => A(9), Z => n35);
   U59 : NAND3_X1 port map( A1 => n36, A2 => n85, A3 => n35, ZN => p(10));
   U60 : MUX2_X1 port map( A => n90, B => n70, S => A(11), Z => n39);
   U61 : MUX2_X1 port map( A => n5, B => n87, S => A(10), Z => n38);
   U62 : NAND3_X1 port map( A1 => n39, A2 => n85, A3 => n38, ZN => p(11));
   U63 : MUX2_X1 port map( A => n88, B => n87, S => A(11), Z => n41);
   U64 : MUX2_X1 port map( A => n92, B => n83, S => A(12), Z => n40);
   U65 : NAND3_X1 port map( A1 => n41, A2 => n85, A3 => n40, ZN => p(12));
   U66 : MUX2_X1 port map( A => n5, B => n87, S => A(12), Z => n43);
   U67 : MUX2_X1 port map( A => n90, B => n70, S => A(13), Z => n42);
   U68 : NAND3_X1 port map( A1 => n43, A2 => n85, A3 => n42, ZN => p(13));
   U69 : NAND3_X1 port map( A1 => b(2), A2 => n45, A3 => n44, ZN => n77);
   U70 : MUX2_X1 port map( A => n77, B => n87, S => A(13), Z => n47);
   U71 : MUX2_X1 port map( A => n4, B => n83, S => A(14), Z => n46);
   U72 : NAND3_X1 port map( A1 => n47, A2 => n85, A3 => n46, ZN => p(14));
   U73 : MUX2_X1 port map( A => n88, B => n87, S => A(14), Z => n49);
   U74 : MUX2_X1 port map( A => n4, B => n6, S => A(15), Z => n48);
   U75 : NAND3_X1 port map( A1 => n49, A2 => n85, A3 => n48, ZN => p(15));
   U76 : MUX2_X1 port map( A => n5, B => n87, S => A(15), Z => n51);
   U77 : MUX2_X1 port map( A => n4, B => n70, S => A(16), Z => n50);
   U78 : NAND3_X1 port map( A1 => n51, A2 => n85, A3 => n50, ZN => p(16));
   U79 : MUX2_X1 port map( A => n77, B => n87, S => A(16), Z => n53);
   U80 : MUX2_X1 port map( A => n4, B => n6, S => A(17), Z => n52);
   U81 : NAND3_X1 port map( A1 => n53, A2 => n85, A3 => n52, ZN => p(17));
   U82 : MUX2_X1 port map( A => n92, B => n70, S => A(18), Z => n55);
   U83 : MUX2_X1 port map( A => n77, B => n87, S => A(17), Z => n54);
   U84 : NAND3_X1 port map( A1 => n55, A2 => n54, A3 => n85, ZN => p(18));
   U85 : MUX2_X1 port map( A => n77, B => n87, S => A(18), Z => n57);
   U86 : MUX2_X1 port map( A => n78, B => n83, S => A(19), Z => n56);
   U87 : NAND3_X1 port map( A1 => n56, A2 => n85, A3 => n57, ZN => p(19));
   U88 : MUX2_X1 port map( A => n77, B => n87, S => A(19), Z => n59);
   U89 : MUX2_X1 port map( A => n90, B => n70, S => A(20), Z => n58);
   U90 : NAND3_X1 port map( A1 => n59, A2 => n58, A3 => n85, ZN => p(20));
   U91 : MUX2_X1 port map( A => n77, B => n87, S => A(20), Z => n61);
   U92 : MUX2_X1 port map( A => n90, B => n83, S => A(21), Z => n60);
   U93 : NAND3_X1 port map( A1 => n61, A2 => n85, A3 => n60, ZN => p(21));
   U94 : MUX2_X1 port map( A => n77, B => n87, S => A(21), Z => n63);
   U95 : MUX2_X1 port map( A => n78, B => n70, S => A(22), Z => n62);
   U96 : NAND3_X1 port map( A1 => n63, A2 => n85, A3 => n62, ZN => p(22));
   U97 : MUX2_X1 port map( A => n77, B => n87, S => A(22), Z => n65);
   U98 : MUX2_X1 port map( A => n90, B => n70, S => A(23), Z => n64);
   U99 : NAND3_X1 port map( A1 => n65, A2 => n85, A3 => n64, ZN => p(23));
   U100 : MUX2_X1 port map( A => n88, B => n87, S => A(23), Z => n67);
   U101 : MUX2_X1 port map( A => n78, B => n83, S => n93, Z => n66);
   U102 : NAND3_X1 port map( A1 => n67, A2 => n85, A3 => n66, ZN => p(24));
   U103 : MUX2_X1 port map( A => n78, B => n70, S => n93, Z => n69);
   U104 : MUX2_X1 port map( A => n77, B => n87, S => n93, Z => n68);
   U105 : NAND3_X1 port map( A1 => n85, A2 => n69, A3 => n68, ZN => p(25));
   U106 : MUX2_X1 port map( A => n5, B => n87, S => n93, Z => n72);
   U107 : MUX2_X1 port map( A => n90, B => n70, S => n93, Z => n71);
   U108 : NAND3_X1 port map( A1 => n72, A2 => n85, A3 => n71, ZN => p(26));
   U109 : MUX2_X1 port map( A => n77, B => n87, S => n93, Z => n74);
   U110 : MUX2_X1 port map( A => n4, B => n6, S => n93, Z => n73);
   U111 : NAND3_X1 port map( A1 => n74, A2 => n85, A3 => n73, ZN => p(27));
   U112 : MUX2_X1 port map( A => n88, B => n87, S => n93, Z => n76);
   U113 : MUX2_X1 port map( A => n90, B => n6, S => n93, Z => n75);
   U114 : NAND3_X1 port map( A1 => n76, A2 => n85, A3 => n75, ZN => p(28));
   U115 : MUX2_X1 port map( A => n77, B => n87, S => n93, Z => n80);
   U116 : MUX2_X1 port map( A => n78, B => n83, S => n93, Z => n79);
   U117 : NAND3_X1 port map( A1 => n80, A2 => n85, A3 => n79, ZN => p(29));
   U118 : MUX2_X1 port map( A => n5, B => n87, S => n93, Z => n82);
   U119 : MUX2_X1 port map( A => n92, B => n6, S => n93, Z => n81);
   U120 : NAND3_X1 port map( A1 => n82, A2 => n85, A3 => n81, ZN => p(30));
   U121 : MUX2_X1 port map( A => n88, B => n87, S => n93, Z => n86);
   U122 : MUX2_X1 port map( A => n4, B => n6, S => n93, Z => n84);
   U123 : NAND3_X1 port map( A1 => n86, A2 => n85, A3 => n84, ZN => p(31));
   U124 : MUX2_X1 port map( A => n5, B => n87, S => n93, Z => n89);
   U125 : NAND2_X1 port map( A1 => n4, A2 => n89, ZN => p(32));
   U21 : INV_X1 port map( A => b(2), ZN => n37);
   U18 : INV_X1 port map( A => b(1), ZN => n44);
   U10 : NAND2_X1 port map( A1 => n13, A2 => n37, ZN => n6);
   U12 : NAND2_X1 port map( A1 => b(2), A2 => n24, ZN => n92);
   n93 <= '0';
   U5 : NAND2_X2 port map( A1 => b(0), A2 => b(1), ZN => n87);
   U6 : NAND3_X2 port map( A1 => b(0), A2 => b(1), A3 => b(2), ZN => n85);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_12 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_12;

architecture SYN_beh of ENC_12 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net32441, net32448, net32450, net32452, net32457, net32474, net32475,
      net32478, net32479, net32518, net32519, net32520, net33933, net32480, 
      net32453, net32446, n2, n3, n4, n7, n8, n9, n10, n12, n13, n14, n15, n16,
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71 : std_logic;

begin
   
   U4 : NAND2_X1 port map( A1 => n7, A2 => n2, ZN => n3);
   U5 : NAND2_X1 port map( A1 => net32519, A2 => A(20), ZN => n4);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n52);
   U7 : INV_X1 port map( A => A(20), ZN => n2);
   U16 : MUX2_X1 port map( A => n7, B => net32519, S => n71, Z => n8);
   U17 : NAND3_X1 port map( A1 => net32453, A2 => net32446, A3 => n8, ZN => 
                           p(29));
   U20 : MUX2_X1 port map( A => net32441, B => n12, S => n71, Z => net32457);
   U25 : XNOR2_X1 port map( A => b(0), B => n10, ZN => net33933);
   U26 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => net32480);
   U27 : INV_X1 port map( A => b(0), ZN => n9);
   U28 : XOR2_X1 port map( A => b(1), B => b(0), Z => net32478);
   U30 : NAND3_X1 port map( A1 => net32474, A2 => net32446, A3 => net32475, ZN 
                           => p(19));
   U32 : MUX2_X1 port map( A => net32448, B => net32452, S => n71, Z => 
                           net32453);
   U38 : MUX2_X1 port map( A => n7, B => net32519, S => n71, Z => net32450);
   U39 : MUX2_X1 port map( A => net32518, B => net32452, S => A(0), Z => 
                           net32520);
   U40 : NAND2_X1 port map( A1 => net32480, A2 => b(2), ZN => net32441);
   U43 : NAND2_X1 port map( A1 => net33933, A2 => net32479, ZN => n12);
   U49 : NAND2_X1 port map( A1 => b(2), A2 => net32519, ZN => net32518);
   U50 : OAI211_X1 port map( C1 => net32479, C2 => net32519, A => n7, B => 
                           net32520, ZN => p(0));
   U51 : MUX2_X1 port map( A => n7, B => net32519, S => A(0), Z => n14);
   U52 : MUX2_X1 port map( A => net32448, B => net32452, S => A(1), Z => n13);
   U53 : NAND3_X1 port map( A1 => n14, A2 => net32446, A3 => n13, ZN => p(1));
   U54 : MUX2_X1 port map( A => n7, B => net32519, S => A(1), Z => n16);
   U55 : MUX2_X1 port map( A => net32448, B => net32452, S => A(2), Z => n15);
   U56 : NAND3_X1 port map( A1 => n16, A2 => net32446, A3 => n15, ZN => p(2));
   U57 : MUX2_X1 port map( A => n7, B => net32519, S => A(2), Z => n18);
   U58 : MUX2_X1 port map( A => net32441, B => n12, S => A(3), Z => n17);
   U59 : NAND3_X1 port map( A1 => n18, A2 => net32446, A3 => n17, ZN => p(3));
   U60 : MUX2_X1 port map( A => n7, B => net32519, S => A(3), Z => n20);
   U61 : MUX2_X1 port map( A => net32448, B => net32452, S => A(4), Z => n19);
   U62 : NAND3_X1 port map( A1 => n20, A2 => net32446, A3 => n19, ZN => p(4));
   U63 : MUX2_X1 port map( A => n7, B => net32519, S => A(4), Z => n22);
   U64 : MUX2_X1 port map( A => net32441, B => net32452, S => A(5), Z => n21);
   U65 : NAND3_X1 port map( A1 => n22, A2 => net32446, A3 => n21, ZN => p(5));
   U66 : MUX2_X1 port map( A => n7, B => net32519, S => A(5), Z => n24);
   U67 : MUX2_X1 port map( A => net32448, B => net32452, S => A(6), Z => n23);
   U68 : NAND3_X1 port map( A1 => n24, A2 => net32446, A3 => n23, ZN => p(6));
   U69 : MUX2_X1 port map( A => n7, B => net32519, S => A(6), Z => n26);
   U70 : MUX2_X1 port map( A => net32448, B => net32452, S => A(7), Z => n25);
   U71 : NAND3_X1 port map( A1 => n26, A2 => net32446, A3 => n25, ZN => p(7));
   U72 : MUX2_X1 port map( A => n7, B => net32519, S => A(7), Z => n28);
   U73 : MUX2_X1 port map( A => net32441, B => net32452, S => A(8), Z => n27);
   U74 : NAND3_X1 port map( A1 => n28, A2 => net32446, A3 => n27, ZN => p(8));
   U75 : MUX2_X1 port map( A => n7, B => net32519, S => A(8), Z => n30);
   U76 : MUX2_X1 port map( A => net32441, B => net32452, S => A(9), Z => n29);
   U77 : NAND3_X1 port map( A1 => n30, A2 => net32446, A3 => n29, ZN => p(9));
   U78 : MUX2_X1 port map( A => n7, B => net32519, S => A(9), Z => n32);
   U79 : MUX2_X1 port map( A => net32441, B => net32452, S => A(10), Z => n31);
   U80 : NAND3_X1 port map( A1 => n32, A2 => net32446, A3 => n31, ZN => p(10));
   U81 : MUX2_X1 port map( A => n7, B => net32519, S => A(10), Z => n34);
   U82 : MUX2_X1 port map( A => net32448, B => net32452, S => A(11), Z => n33);
   U83 : NAND3_X1 port map( A1 => n34, A2 => net32446, A3 => n33, ZN => p(11));
   U84 : MUX2_X1 port map( A => n7, B => net32519, S => A(11), Z => n36);
   U85 : MUX2_X1 port map( A => net32441, B => net32452, S => A(12), Z => n35);
   U86 : NAND3_X1 port map( A1 => n36, A2 => net32446, A3 => n35, ZN => p(12));
   U87 : MUX2_X1 port map( A => n7, B => net32519, S => A(12), Z => n38);
   U88 : MUX2_X1 port map( A => net32441, B => net32452, S => A(13), Z => n37);
   U89 : NAND3_X1 port map( A1 => n38, A2 => net32446, A3 => n37, ZN => p(13));
   U90 : MUX2_X1 port map( A => net32448, B => n12, S => A(14), Z => n40);
   U91 : MUX2_X1 port map( A => n7, B => net32519, S => A(13), Z => n39);
   U92 : NAND3_X1 port map( A1 => n40, A2 => net32446, A3 => n39, ZN => p(14));
   U93 : MUX2_X1 port map( A => n7, B => net32519, S => A(14), Z => n42);
   U94 : MUX2_X1 port map( A => net32448, B => net32452, S => A(15), Z => n41);
   U95 : NAND3_X1 port map( A1 => n42, A2 => net32446, A3 => n41, ZN => p(15));
   U96 : MUX2_X1 port map( A => n7, B => net32519, S => A(15), Z => n44);
   U97 : MUX2_X1 port map( A => net32448, B => n12, S => A(16), Z => n43);
   U98 : NAND3_X1 port map( A1 => n44, A2 => net32446, A3 => n43, ZN => p(16));
   U99 : MUX2_X1 port map( A => n7, B => net32519, S => A(16), Z => n46);
   U100 : MUX2_X1 port map( A => net32441, B => net32452, S => A(17), Z => n45)
                           ;
   U101 : NAND3_X1 port map( A1 => n46, A2 => net32446, A3 => n45, ZN => p(17))
                           ;
   U102 : NAND2_X1 port map( A1 => net32478, A2 => net32479, ZN => n67);
   U103 : MUX2_X1 port map( A => net32448, B => n67, S => A(18), Z => n48);
   U104 : MUX2_X1 port map( A => n7, B => net32519, S => A(17), Z => n47);
   U105 : NAND3_X1 port map( A1 => n48, A2 => net32446, A3 => n47, ZN => p(18))
                           ;
   U106 : MUX2_X1 port map( A => n7, B => net32519, S => A(18), Z => net32474);
   U107 : MUX2_X1 port map( A => net32448, B => n12, S => A(19), Z => net32475)
                           ;
   U108 : MUX2_X1 port map( A => n7, B => net32519, S => A(19), Z => n50);
   U109 : MUX2_X1 port map( A => net32448, B => n12, S => A(20), Z => n49);
   U110 : NAND3_X1 port map( A1 => n50, A2 => net32446, A3 => n49, ZN => p(20))
                           ;
   U111 : MUX2_X1 port map( A => net32441, B => n12, S => A(21), Z => n51);
   U112 : NAND3_X1 port map( A1 => n52, A2 => net32446, A3 => n51, ZN => p(21))
                           ;
   U113 : MUX2_X1 port map( A => n7, B => net32519, S => A(21), Z => n54);
   U114 : MUX2_X1 port map( A => net32441, B => net32452, S => A(22), Z => n53)
                           ;
   U115 : NAND3_X1 port map( A1 => n54, A2 => net32446, A3 => n53, ZN => p(22))
                           ;
   U116 : MUX2_X1 port map( A => n7, B => net32519, S => A(22), Z => n56);
   U117 : MUX2_X1 port map( A => net32441, B => net32452, S => A(23), Z => n55)
                           ;
   U118 : NAND3_X1 port map( A1 => n56, A2 => net32446, A3 => n55, ZN => p(23))
                           ;
   U119 : MUX2_X1 port map( A => n7, B => net32519, S => A(23), Z => n58);
   U120 : MUX2_X1 port map( A => net32441, B => net32452, S => n71, Z => n57);
   U121 : NAND3_X1 port map( A1 => n58, A2 => net32446, A3 => n57, ZN => p(24))
                           ;
   U122 : MUX2_X1 port map( A => n7, B => net32519, S => n71, Z => n60);
   U123 : MUX2_X1 port map( A => net32441, B => net32452, S => n71, Z => n59);
   U124 : NAND3_X1 port map( A1 => n60, A2 => net32446, A3 => n59, ZN => p(25))
                           ;
   U125 : MUX2_X1 port map( A => net32448, B => net32452, S => n71, Z => n62);
   U126 : MUX2_X1 port map( A => n7, B => net32519, S => n71, Z => n61);
   U127 : NAND3_X1 port map( A1 => n62, A2 => net32446, A3 => n61, ZN => p(26))
                           ;
   U128 : MUX2_X1 port map( A => net32448, B => n12, S => n71, Z => n64);
   U129 : MUX2_X1 port map( A => n7, B => net32519, S => n71, Z => n63);
   U130 : NAND3_X1 port map( A1 => net32446, A2 => n64, A3 => n63, ZN => p(27))
                           ;
   U131 : MUX2_X1 port map( A => n7, B => net32519, S => n71, Z => n65);
   U132 : NAND3_X1 port map( A1 => n65, A2 => net32446, A3 => net32457, ZN => 
                           p(28));
   U133 : MUX2_X1 port map( A => net32441, B => n12, S => n71, Z => n66);
   U134 : NAND3_X1 port map( A1 => net32450, A2 => n66, A3 => net32446, ZN => 
                           p(30));
   U135 : MUX2_X1 port map( A => n7, B => net32519, S => n71, Z => n69);
   U136 : MUX2_X1 port map( A => net32448, B => n67, S => n71, Z => n68);
   U137 : NAND3_X1 port map( A1 => n69, A2 => net32446, A3 => n68, ZN => p(31))
                           ;
   U138 : MUX2_X1 port map( A => n7, B => net32519, S => n71, Z => n70);
   U139 : NAND2_X1 port map( A1 => net32441, A2 => n70, ZN => p(32));
   U36 : INV_X1 port map( A => b(2), ZN => net32479);
   U21 : NAND2_X2 port map( A1 => b(0), A2 => b(1), ZN => net32519);
   U24 : INV_X1 port map( A => b(1), ZN => n10);
   U22 : NAND3_X2 port map( A1 => n9, A2 => b(2), A3 => n10, ZN => n7);
   U35 : NAND2_X1 port map( A1 => net33933, A2 => net32479, ZN => net32452);
   U8 : NAND2_X1 port map( A1 => net32480, A2 => b(2), ZN => net32448);
   n71 <= '0';
   U3 : NAND2_X2 port map( A1 => b(2), A2 => net32518, ZN => net32446);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_13 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_13;

architecture SYN_beh of ENC_13 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n11, n12, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, 
      n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47
      , n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, 
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n104 : 
      std_logic;

begin
   
   U5 : NAND2_X1 port map( A1 => n56, A2 => n63, ZN => n1);
   U9 : OR2_X1 port map( A1 => n23, A2 => b(2), ZN => n12);
   U13 : NAND2_X1 port map( A1 => n49, A2 => n95, ZN => n5);
   U25 : XNOR2_X1 port map( A => n63, B => b(0), ZN => n11);
   U26 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n23);
   U27 : NAND3_X1 port map( A1 => b(0), A2 => b(1), A3 => b(2), ZN => n25);
   U29 : INV_X1 port map( A => b(0), ZN => n56);
   U32 : MUX2_X1 port map( A => n95, B => n12, S => A(0), Z => n24);
   U33 : NAND3_X1 port map( A1 => n25, A2 => n94, A3 => n24, ZN => p(0));
   U35 : MUX2_X1 port map( A => n94, B => n99, S => A(0), Z => n27);
   U37 : NAND2_X1 port map( A1 => n56, A2 => n63, ZN => n48);
   U39 : MUX2_X1 port map( A => n102, B => n91, S => A(1), Z => n26);
   U40 : NAND3_X1 port map( A1 => n27, A2 => n97, A3 => n26, ZN => p(1));
   U41 : MUX2_X1 port map( A => n94, B => n99, S => A(1), Z => n29);
   U42 : MUX2_X1 port map( A => n102, B => n12, S => A(2), Z => n28);
   U43 : NAND3_X1 port map( A1 => n29, A2 => n97, A3 => n28, ZN => p(2));
   U44 : MUX2_X1 port map( A => n94, B => n99, S => A(2), Z => n31);
   U45 : MUX2_X1 port map( A => n102, B => n91, S => A(3), Z => n30);
   U46 : NAND3_X1 port map( A1 => n31, A2 => n97, A3 => n30, ZN => p(3));
   U47 : MUX2_X1 port map( A => n94, B => n99, S => A(3), Z => n33);
   U48 : MUX2_X1 port map( A => n79, B => n12, S => A(4), Z => n32);
   U49 : NAND3_X1 port map( A1 => n33, A2 => n97, A3 => n32, ZN => p(4));
   U50 : MUX2_X1 port map( A => n94, B => n99, S => A(4), Z => n35);
   U51 : MUX2_X1 port map( A => n79, B => n91, S => A(5), Z => n34);
   U52 : NAND3_X1 port map( A1 => n35, A2 => n97, A3 => n34, ZN => p(5));
   U53 : MUX2_X1 port map( A => n94, B => n99, S => A(5), Z => n37);
   U54 : MUX2_X1 port map( A => n79, B => n91, S => A(6), Z => n36);
   U55 : NAND3_X1 port map( A1 => n37, A2 => n97, A3 => n36, ZN => p(6));
   U56 : MUX2_X1 port map( A => n94, B => n99, S => A(6), Z => n39);
   U57 : MUX2_X1 port map( A => n102, B => n91, S => A(7), Z => n38);
   U58 : NAND3_X1 port map( A1 => n39, A2 => n97, A3 => n38, ZN => p(7));
   U59 : MUX2_X1 port map( A => n94, B => n99, S => A(7), Z => n41);
   U60 : MUX2_X1 port map( A => n102, B => n12, S => A(8), Z => n40);
   U61 : NAND3_X1 port map( A1 => n41, A2 => n97, A3 => n40, ZN => p(8));
   U62 : MUX2_X1 port map( A => n94, B => n99, S => A(8), Z => n43);
   U63 : MUX2_X1 port map( A => n102, B => n12, S => A(9), Z => n42);
   U64 : NAND3_X1 port map( A1 => n43, A2 => n97, A3 => n42, ZN => p(9));
   U65 : MUX2_X1 port map( A => n94, B => n99, S => A(9), Z => n45);
   U66 : MUX2_X1 port map( A => n102, B => n91, S => A(10), Z => n44);
   U67 : NAND3_X1 port map( A1 => n45, A2 => n97, A3 => n44, ZN => p(10));
   U68 : MUX2_X1 port map( A => n94, B => n99, S => A(10), Z => n47);
   U69 : MUX2_X1 port map( A => n102, B => n91, S => A(11), Z => n46);
   U70 : NAND3_X1 port map( A1 => n47, A2 => n97, A3 => n46, ZN => p(11));
   U72 : XOR2_X1 port map( A => b(0), B => b(1), Z => n49);
   U73 : NAND2_X1 port map( A1 => n49, A2 => n95, ZN => n88);
   U74 : MUX2_X1 port map( A => n79, B => n88, S => A(12), Z => n51);
   U75 : MUX2_X1 port map( A => n94, B => n99, S => A(11), Z => n50);
   U76 : NAND3_X1 port map( A1 => n51, A2 => n97, A3 => n50, ZN => p(12));
   U77 : MUX2_X1 port map( A => n94, B => n99, S => A(12), Z => n53);
   U78 : MUX2_X1 port map( A => n102, B => n91, S => A(13), Z => n52);
   U79 : NAND3_X1 port map( A1 => n53, A2 => n97, A3 => n52, ZN => p(13));
   U80 : MUX2_X1 port map( A => n94, B => n99, S => A(13), Z => n55);
   U81 : MUX2_X1 port map( A => n102, B => n91, S => A(14), Z => n54);
   U82 : NAND3_X1 port map( A1 => n55, A2 => n97, A3 => n54, ZN => p(14));
   U83 : NAND3_X1 port map( A1 => b(2), A2 => n56, A3 => n63, ZN => n100);
   U84 : MUX2_X1 port map( A => n100, B => n99, S => A(14), Z => n58);
   U85 : MUX2_X1 port map( A => n102, B => n5, S => A(15), Z => n57);
   U86 : NAND3_X1 port map( A1 => n58, A2 => n97, A3 => n57, ZN => p(15));
   U87 : MUX2_X1 port map( A => n100, B => n99, S => A(15), Z => n60);
   U88 : MUX2_X1 port map( A => n102, B => n91, S => A(16), Z => n59);
   U89 : NAND3_X1 port map( A1 => n59, A2 => n97, A3 => n60, ZN => p(16));
   U90 : MUX2_X1 port map( A => n94, B => n99, S => A(16), Z => n62);
   U91 : MUX2_X1 port map( A => n79, B => n91, S => A(17), Z => n61);
   U92 : NAND3_X1 port map( A1 => n62, A2 => n97, A3 => n61, ZN => p(17));
   U93 : NAND2_X1 port map( A1 => n11, A2 => n95, ZN => n64);
   U94 : MUX2_X1 port map( A => n79, B => n64, S => A(18), Z => n66);
   U95 : MUX2_X1 port map( A => n100, B => n99, S => A(17), Z => n65);
   U96 : NAND3_X1 port map( A1 => n66, A2 => n97, A3 => n65, ZN => p(18));
   U97 : MUX2_X1 port map( A => n94, B => n99, S => A(18), Z => n68);
   U98 : MUX2_X1 port map( A => n102, B => n91, S => A(19), Z => n67);
   U99 : NAND3_X1 port map( A1 => n68, A2 => n97, A3 => n67, ZN => p(19));
   U100 : MUX2_X1 port map( A => n100, B => n99, S => A(19), Z => n70);
   U101 : MUX2_X1 port map( A => n79, B => n91, S => A(20), Z => n69);
   U102 : NAND3_X1 port map( A1 => n69, A2 => n70, A3 => n97, ZN => p(20));
   U103 : MUX2_X1 port map( A => n100, B => n99, S => A(20), Z => n72);
   U104 : MUX2_X1 port map( A => n79, B => n5, S => A(21), Z => n71);
   U105 : NAND3_X1 port map( A1 => n72, A2 => n97, A3 => n71, ZN => p(21));
   U106 : MUX2_X1 port map( A => n102, B => n88, S => A(22), Z => n74);
   U107 : MUX2_X1 port map( A => n94, B => n99, S => A(21), Z => n73);
   U108 : NAND3_X1 port map( A1 => n74, A2 => n97, A3 => n73, ZN => p(22));
   U109 : MUX2_X1 port map( A => n79, B => n12, S => A(23), Z => n76);
   U110 : MUX2_X1 port map( A => n94, B => n99, S => A(22), Z => n75);
   U111 : NAND3_X1 port map( A1 => n97, A2 => n76, A3 => n75, ZN => p(23));
   U112 : MUX2_X1 port map( A => n79, B => n5, S => n104, Z => n78);
   U113 : MUX2_X1 port map( A => n100, B => n99, S => A(23), Z => n77);
   U114 : NAND3_X1 port map( A1 => n78, A2 => n97, A3 => n77, ZN => p(24));
   U115 : MUX2_X1 port map( A => n100, B => n99, S => n104, Z => n81);
   U116 : MUX2_X1 port map( A => n79, B => n5, S => n104, Z => n80);
   U117 : NAND3_X1 port map( A1 => n81, A2 => n97, A3 => n80, ZN => p(25));
   U118 : MUX2_X1 port map( A => n100, B => n99, S => n104, Z => n83);
   U119 : MUX2_X1 port map( A => n102, B => n88, S => n104, Z => n82);
   U120 : NAND3_X1 port map( A1 => n83, A2 => n97, A3 => n82, ZN => p(26));
   U121 : MUX2_X1 port map( A => n94, B => n99, S => n104, Z => n85);
   U122 : MUX2_X1 port map( A => n102, B => n91, S => n104, Z => n84);
   U123 : NAND3_X1 port map( A1 => n85, A2 => n97, A3 => n84, ZN => p(27));
   U124 : MUX2_X1 port map( A => n94, B => n99, S => n104, Z => n87);
   U125 : MUX2_X1 port map( A => n102, B => n91, S => n104, Z => n86);
   U126 : NAND3_X1 port map( A1 => n87, A2 => n97, A3 => n86, ZN => p(28));
   U127 : MUX2_X1 port map( A => n94, B => n99, S => n104, Z => n90);
   U128 : MUX2_X1 port map( A => n79, B => n88, S => n104, Z => n89);
   U129 : NAND3_X1 port map( A1 => n90, A2 => n97, A3 => n89, ZN => p(29));
   U130 : MUX2_X1 port map( A => n94, B => n99, S => n104, Z => n93);
   U131 : MUX2_X1 port map( A => n79, B => n12, S => n104, Z => n92);
   U132 : NAND3_X1 port map( A1 => n93, A2 => n97, A3 => n92, ZN => p(30));
   U133 : MUX2_X1 port map( A => n94, B => n99, S => n104, Z => n98);
   U134 : MUX2_X1 port map( A => n102, B => n64, S => n104, Z => n96);
   U135 : NAND3_X1 port map( A1 => n98, A2 => n97, A3 => n96, ZN => p(31));
   U136 : MUX2_X1 port map( A => n100, B => n99, S => n104, Z => n101);
   U137 : NAND2_X1 port map( A1 => n79, A2 => n101, ZN => p(32));
   U31 : INV_X1 port map( A => b(2), ZN => n95);
   U71 : NAND2_X1 port map( A1 => n1, A2 => b(2), ZN => n79);
   U30 : NAND3_X1 port map( A1 => n56, A2 => n63, A3 => b(2), ZN => n94);
   U38 : NAND2_X1 port map( A1 => n48, A2 => b(2), ZN => n102);
   U4 : NAND3_X2 port map( A1 => b(1), A2 => b(2), A3 => b(0), ZN => n97);
   U7 : OR2_X1 port map( A1 => n23, A2 => b(2), ZN => n91);
   U8 : INV_X1 port map( A => b(1), ZN => n63);
   n104 <= '0';
   U3 : NAND2_X2 port map( A1 => b(0), A2 => b(1), ZN => n99);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_14 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_14;

architecture SYN_beh of ENC_14 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43
      , n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, 
      n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72
      , n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n94, n96 : std_logic;

begin
   
   U4 : XNOR2_X1 port map( A => b(0), B => n17, ZN => n18);
   U5 : XNOR2_X1 port map( A => b(0), B => n17, ZN => n48);
   U12 : NAND2_X1 port map( A1 => n18, A2 => n47, ZN => n81);
   U20 : NAND2_X1 port map( A1 => n94, A2 => n90, ZN => p(32));
   U23 : NAND3_X1 port map( A1 => b(0), A2 => b(1), A3 => b(2), ZN => n20);
   U28 : MUX2_X1 port map( A => n47, B => n81, S => A(0), Z => n19);
   U29 : NAND3_X1 port map( A1 => n20, A2 => n89, A3 => n19, ZN => p(0));
   U31 : MUX2_X1 port map( A => n89, B => n88, S => A(0), Z => n22);
   U33 : OAI21_X1 port map( B1 => b(0), B2 => b(1), A => b(2), ZN => n91);
   U34 : MUX2_X1 port map( A => n94, B => n6, S => A(1), Z => n21);
   U35 : NAND3_X1 port map( A1 => n22, A2 => n86, A3 => n21, ZN => p(1));
   U36 : MUX2_X1 port map( A => n89, B => n88, S => A(1), Z => n24);
   U37 : MUX2_X1 port map( A => n91, B => n6, S => A(2), Z => n23);
   U38 : NAND3_X1 port map( A1 => n24, A2 => n86, A3 => n23, ZN => p(2));
   U39 : MUX2_X1 port map( A => n89, B => n88, S => A(2), Z => n26);
   U40 : MUX2_X1 port map( A => n94, B => n6, S => A(3), Z => n25);
   U41 : NAND3_X1 port map( A1 => n26, A2 => n86, A3 => n25, ZN => p(3));
   U42 : MUX2_X1 port map( A => n89, B => n88, S => A(3), Z => n28);
   U43 : MUX2_X1 port map( A => n91, B => n81, S => A(4), Z => n27);
   U44 : NAND3_X1 port map( A1 => n28, A2 => n86, A3 => n27, ZN => p(4));
   U45 : MUX2_X1 port map( A => n89, B => n88, S => A(4), Z => n30);
   U46 : MUX2_X1 port map( A => n94, B => n6, S => A(5), Z => n29);
   U47 : NAND3_X1 port map( A1 => n30, A2 => n86, A3 => n29, ZN => p(5));
   U48 : MUX2_X1 port map( A => n89, B => n88, S => A(5), Z => n32);
   U49 : MUX2_X1 port map( A => n94, B => n6, S => A(6), Z => n31);
   U50 : NAND3_X1 port map( A1 => n32, A2 => n86, A3 => n31, ZN => p(6));
   U51 : MUX2_X1 port map( A => n89, B => n88, S => A(6), Z => n34);
   U52 : MUX2_X1 port map( A => n94, B => n6, S => A(7), Z => n33);
   U53 : NAND3_X1 port map( A1 => n34, A2 => n86, A3 => n33, ZN => p(7));
   U54 : MUX2_X1 port map( A => n89, B => n88, S => A(7), Z => n36);
   U55 : MUX2_X1 port map( A => n94, B => n6, S => A(8), Z => n35);
   U56 : NAND3_X1 port map( A1 => n36, A2 => n86, A3 => n35, ZN => p(8));
   U57 : MUX2_X1 port map( A => n89, B => n88, S => A(8), Z => n38);
   U58 : MUX2_X1 port map( A => n94, B => n6, S => A(9), Z => n37);
   U59 : NAND3_X1 port map( A1 => n38, A2 => n86, A3 => n37, ZN => p(9));
   U60 : MUX2_X1 port map( A => n89, B => n88, S => A(9), Z => n40);
   U61 : MUX2_X1 port map( A => n91, B => n6, S => A(10), Z => n39);
   U62 : NAND3_X1 port map( A1 => n40, A2 => n86, A3 => n39, ZN => p(10));
   U63 : MUX2_X1 port map( A => n89, B => n88, S => A(10), Z => n42);
   U64 : MUX2_X1 port map( A => n91, B => n81, S => A(11), Z => n41);
   U65 : NAND3_X1 port map( A1 => n42, A2 => n86, A3 => n41, ZN => p(11));
   U66 : MUX2_X1 port map( A => n89, B => n88, S => A(11), Z => n44);
   U67 : MUX2_X1 port map( A => n91, B => n6, S => A(12), Z => n43);
   U68 : NAND3_X1 port map( A1 => n44, A2 => n86, A3 => n43, ZN => p(12));
   U69 : MUX2_X1 port map( A => n89, B => n88, S => A(12), Z => n46);
   U70 : MUX2_X1 port map( A => n94, B => n6, S => A(13), Z => n45);
   U71 : NAND3_X1 port map( A1 => n46, A2 => n86, A3 => n45, ZN => p(13));
   U72 : MUX2_X1 port map( A => n94, B => n84, S => A(14), Z => n50);
   U73 : MUX2_X1 port map( A => n89, B => n88, S => A(13), Z => n49);
   U74 : NAND3_X1 port map( A1 => n50, A2 => n86, A3 => n49, ZN => p(14));
   U75 : MUX2_X1 port map( A => n89, B => n88, S => A(14), Z => n52);
   U76 : MUX2_X1 port map( A => n94, B => n84, S => A(15), Z => n51);
   U77 : NAND3_X1 port map( A1 => n52, A2 => n86, A3 => n51, ZN => p(15));
   U78 : MUX2_X1 port map( A => n89, B => n88, S => A(15), Z => n54);
   U79 : MUX2_X1 port map( A => n94, B => n81, S => A(16), Z => n53);
   U80 : NAND3_X1 port map( A1 => n54, A2 => n86, A3 => n53, ZN => p(16));
   U81 : MUX2_X1 port map( A => n89, B => n88, S => A(16), Z => n56);
   U82 : MUX2_X1 port map( A => n94, B => n84, S => A(17), Z => n55);
   U83 : NAND3_X1 port map( A1 => n56, A2 => n86, A3 => n55, ZN => p(17));
   U84 : MUX2_X1 port map( A => n89, B => n88, S => A(17), Z => n58);
   U85 : MUX2_X1 port map( A => n94, B => n6, S => A(18), Z => n57);
   U86 : NAND3_X1 port map( A1 => n58, A2 => n86, A3 => n57, ZN => p(18));
   U87 : MUX2_X1 port map( A => n89, B => n88, S => A(18), Z => n60);
   U88 : MUX2_X1 port map( A => n94, B => n81, S => A(19), Z => n59);
   U89 : NAND3_X1 port map( A1 => n60, A2 => n86, A3 => n59, ZN => p(19));
   U90 : MUX2_X1 port map( A => n89, B => n88, S => A(19), Z => n62);
   U91 : MUX2_X1 port map( A => n91, B => n84, S => A(20), Z => n61);
   U92 : NAND3_X1 port map( A1 => n62, A2 => n61, A3 => n86, ZN => p(20));
   U93 : MUX2_X1 port map( A => n89, B => n88, S => A(20), Z => n64);
   U94 : MUX2_X1 port map( A => n94, B => n84, S => A(21), Z => n63);
   U95 : NAND3_X1 port map( A1 => n64, A2 => n86, A3 => n63, ZN => p(21));
   U96 : MUX2_X1 port map( A => n89, B => n88, S => A(21), Z => n66);
   U97 : MUX2_X1 port map( A => n94, B => n84, S => A(22), Z => n65);
   U98 : NAND3_X1 port map( A1 => n66, A2 => n86, A3 => n65, ZN => p(22));
   U99 : MUX2_X1 port map( A => n89, B => n88, S => A(22), Z => n68);
   U100 : MUX2_X1 port map( A => n94, B => n84, S => A(23), Z => n67);
   U101 : NAND3_X1 port map( A1 => n68, A2 => n86, A3 => n67, ZN => p(23));
   U102 : MUX2_X1 port map( A => n94, B => n84, S => n96, Z => n70);
   U103 : MUX2_X1 port map( A => n89, B => n88, S => A(23), Z => n69);
   U104 : NAND3_X1 port map( A1 => n70, A2 => n86, A3 => n69, ZN => p(24));
   U105 : MUX2_X1 port map( A => n89, B => n88, S => n96, Z => n72);
   U106 : MUX2_X1 port map( A => n94, B => n84, S => n96, Z => n71);
   U107 : NAND3_X1 port map( A1 => n72, A2 => n86, A3 => n71, ZN => p(25));
   U108 : MUX2_X1 port map( A => n89, B => n88, S => n96, Z => n74);
   U109 : MUX2_X1 port map( A => n91, B => n84, S => n96, Z => n73);
   U110 : NAND3_X1 port map( A1 => n74, A2 => n73, A3 => n86, ZN => p(26));
   U111 : MUX2_X1 port map( A => n89, B => n88, S => n96, Z => n76);
   U112 : MUX2_X1 port map( A => n94, B => n6, S => n96, Z => n75);
   U113 : NAND3_X1 port map( A1 => n76, A2 => n86, A3 => n75, ZN => p(27));
   U114 : MUX2_X1 port map( A => n89, B => n88, S => n96, Z => n78);
   U115 : MUX2_X1 port map( A => n91, B => n84, S => n96, Z => n77);
   U116 : NAND3_X1 port map( A1 => n78, A2 => n86, A3 => n77, ZN => p(28));
   U117 : MUX2_X1 port map( A => n89, B => n88, S => n96, Z => n80);
   U118 : MUX2_X1 port map( A => n91, B => n84, S => n96, Z => n79);
   U119 : NAND3_X1 port map( A1 => n80, A2 => n86, A3 => n79, ZN => p(29));
   U120 : MUX2_X1 port map( A => n89, B => n88, S => n96, Z => n83);
   U121 : MUX2_X1 port map( A => n94, B => n6, S => n96, Z => n82);
   U122 : NAND3_X1 port map( A1 => n83, A2 => n86, A3 => n82, ZN => p(30));
   U123 : MUX2_X1 port map( A => n89, B => n88, S => n96, Z => n87);
   U124 : MUX2_X1 port map( A => n94, B => n84, S => n96, Z => n85);
   U125 : NAND3_X1 port map( A1 => n87, A2 => n86, A3 => n85, ZN => p(31));
   U126 : MUX2_X1 port map( A => n89, B => n88, S => n96, Z => n90);
   U13 : NAND2_X1 port map( A1 => n48, A2 => n47, ZN => n84);
   U3 : NAND2_X1 port map( A1 => n18, A2 => n47, ZN => n6);
   U26 : NAND3_X2 port map( A1 => n17, A2 => n16, A3 => b(2), ZN => n89);
   U7 : BUF_X2 port map( A => n91, Z => n94);
   U9 : NAND3_X2 port map( A1 => b(1), A2 => b(2), A3 => b(0), ZN => n86);
   U10 : INV_X1 port map( A => b(1), ZN => n17);
   U11 : INV_X1 port map( A => b(2), ZN => n47);
   U14 : INV_X1 port map( A => b(0), ZN => n16);
   n96 <= '0';
   U6 : NAND2_X2 port map( A1 => b(0), A2 => b(1), ZN => n88);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_15 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_15;

architecture SYN_beh of ENC_15 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, 
      n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45, n46, n47, n49, n50, n51, n52, n53, n54, n55, n56, 
      n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71
      , n72, n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, 
      n87, n88, n89, n90, n91, n92, n93, n94, n96, n98, n99 : std_logic;

begin
   
   U4 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n74);
   U12 : NAND2_X1 port map( A1 => n96, A2 => n71, ZN => n83);
   U19 : AND2_X1 port map( A1 => b(2), A2 => n18, ZN => n3);
   U20 : AOI22_X1 port map( A1 => b(2), A2 => n74, B1 => n73, B2 => n99, ZN => 
                           n76);
   U21 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n72);
   U22 : NOR2_X1 port map( A1 => n72, A2 => b(2), ZN => n73);
   U25 : INV_X1 port map( A => b(0), ZN => n18);
   U27 : NAND2_X1 port map( A1 => n3, A2 => n47, ZN => n92);
   U29 : NAND2_X1 port map( A1 => n96, A2 => n71, ZN => n88);
   U30 : MUX2_X1 port map( A => n71, B => n4, S => A(0), Z => n15);
   U31 : OAI211_X1 port map( C1 => n71, C2 => n16, A => n92, B => n15, ZN => 
                           p(0));
   U32 : MUX2_X1 port map( A => n92, B => n16, S => A(0), Z => n20);
   U33 : INV_X1 port map( A => n16, ZN => n17);
   U36 : MUX2_X1 port map( A => n94, B => n88, S => A(1), Z => n19);
   U37 : NAND3_X1 port map( A1 => n20, A2 => n90, A3 => n19, ZN => p(1));
   U38 : MUX2_X1 port map( A => n92, B => n16, S => A(1), Z => n22);
   U39 : MUX2_X1 port map( A => n94, B => n4, S => A(2), Z => n21);
   U40 : NAND3_X1 port map( A1 => n22, A2 => n90, A3 => n21, ZN => p(2));
   U41 : MUX2_X1 port map( A => n92, B => n16, S => A(2), Z => n24);
   U42 : MUX2_X1 port map( A => n94, B => n88, S => A(3), Z => n23);
   U43 : NAND3_X1 port map( A1 => n24, A2 => n90, A3 => n23, ZN => p(3));
   U44 : MUX2_X1 port map( A => n92, B => n16, S => A(3), Z => n26);
   U45 : MUX2_X1 port map( A => n94, B => n4, S => A(4), Z => n25);
   U46 : NAND3_X1 port map( A1 => n26, A2 => n90, A3 => n25, ZN => p(4));
   U47 : MUX2_X1 port map( A => n92, B => n16, S => A(4), Z => n28);
   U48 : MUX2_X1 port map( A => n94, B => n88, S => A(5), Z => n27);
   U49 : NAND3_X1 port map( A1 => n28, A2 => n90, A3 => n27, ZN => p(5));
   U50 : MUX2_X1 port map( A => n92, B => n16, S => A(5), Z => n30);
   U51 : MUX2_X1 port map( A => n94, B => n4, S => A(6), Z => n29);
   U52 : NAND3_X1 port map( A1 => n30, A2 => n90, A3 => n29, ZN => p(6));
   U53 : MUX2_X1 port map( A => n92, B => n16, S => A(6), Z => n32);
   U54 : MUX2_X1 port map( A => n94, B => n88, S => A(7), Z => n31);
   U55 : NAND3_X1 port map( A1 => n32, A2 => n90, A3 => n31, ZN => p(7));
   U56 : MUX2_X1 port map( A => n92, B => n16, S => A(7), Z => n34);
   U57 : MUX2_X1 port map( A => n94, B => n4, S => A(8), Z => n33);
   U58 : NAND3_X1 port map( A1 => n34, A2 => n90, A3 => n33, ZN => p(8));
   U59 : MUX2_X1 port map( A => n92, B => n16, S => A(8), Z => n36);
   U60 : MUX2_X1 port map( A => n94, B => n88, S => A(9), Z => n35);
   U61 : NAND3_X1 port map( A1 => n36, A2 => n90, A3 => n35, ZN => p(9));
   U62 : MUX2_X1 port map( A => n92, B => n16, S => A(9), Z => n38);
   U63 : MUX2_X1 port map( A => n94, B => n4, S => A(10), Z => n37);
   U64 : NAND3_X1 port map( A1 => n38, A2 => n90, A3 => n37, ZN => p(10));
   U65 : MUX2_X1 port map( A => n92, B => n16, S => A(10), Z => n40);
   U66 : MUX2_X1 port map( A => n94, B => n88, S => A(11), Z => n39);
   U67 : NAND3_X1 port map( A1 => n40, A2 => n90, A3 => n39, ZN => p(11));
   U68 : MUX2_X1 port map( A => n92, B => n16, S => A(11), Z => n42);
   U69 : MUX2_X1 port map( A => n94, B => n4, S => A(12), Z => n41);
   U70 : NAND3_X1 port map( A1 => n42, A2 => n90, A3 => n41, ZN => p(12));
   U71 : MUX2_X1 port map( A => n92, B => n16, S => A(12), Z => n44);
   U72 : MUX2_X1 port map( A => n94, B => n88, S => A(13), Z => n43);
   U73 : NAND3_X1 port map( A1 => n44, A2 => n90, A3 => n43, ZN => p(13));
   U74 : MUX2_X1 port map( A => n92, B => n16, S => A(13), Z => n46);
   U75 : MUX2_X1 port map( A => n94, B => n4, S => A(14), Z => n45);
   U76 : NAND3_X1 port map( A1 => n46, A2 => n90, A3 => n45, ZN => p(14));
   U77 : NAND2_X1 port map( A1 => n3, A2 => n47, ZN => n80);
   U78 : MUX2_X1 port map( A => n80, B => n16, S => A(14), Z => n50);
   U79 : MUX2_X1 port map( A => n94, B => n83, S => A(15), Z => n49);
   U80 : NAND3_X1 port map( A1 => n50, A2 => n90, A3 => n49, ZN => p(15));
   U81 : MUX2_X1 port map( A => n98, B => n16, S => A(15), Z => n52);
   U82 : MUX2_X1 port map( A => n94, B => n88, S => A(16), Z => n51);
   U83 : NAND3_X1 port map( A1 => n52, A2 => n90, A3 => n51, ZN => p(16));
   U84 : MUX2_X1 port map( A => n98, B => n16, S => A(16), Z => n54);
   U85 : MUX2_X1 port map( A => n94, B => n4, S => A(17), Z => n53);
   U86 : NAND3_X1 port map( A1 => n54, A2 => n90, A3 => n53, ZN => p(17));
   U87 : MUX2_X1 port map( A => n98, B => n16, S => A(17), Z => n56);
   U88 : MUX2_X1 port map( A => n94, B => n88, S => A(18), Z => n55);
   U89 : NAND3_X1 port map( A1 => n56, A2 => n90, A3 => n55, ZN => p(18));
   U90 : MUX2_X1 port map( A => n98, B => n16, S => A(18), Z => n58);
   U91 : MUX2_X1 port map( A => n94, B => n83, S => A(19), Z => n57);
   U92 : NAND3_X1 port map( A1 => n58, A2 => n90, A3 => n57, ZN => p(19));
   U93 : MUX2_X1 port map( A => n98, B => n16, S => A(19), Z => n60);
   U94 : MUX2_X1 port map( A => n94, B => n4, S => A(20), Z => n59);
   U95 : NAND3_X1 port map( A1 => n60, A2 => n90, A3 => n59, ZN => p(20));
   U96 : MUX2_X1 port map( A => n98, B => n16, S => A(20), Z => n62);
   U97 : MUX2_X1 port map( A => n94, B => n83, S => A(21), Z => n61);
   U98 : NAND3_X1 port map( A1 => n62, A2 => n90, A3 => n61, ZN => p(21));
   U99 : MUX2_X1 port map( A => n80, B => n16, S => A(21), Z => n64);
   U100 : MUX2_X1 port map( A => n94, B => n83, S => A(22), Z => n63);
   U101 : NAND3_X1 port map( A1 => n64, A2 => n90, A3 => n63, ZN => p(22));
   U102 : MUX2_X1 port map( A => n80, B => n16, S => A(22), Z => n66);
   U103 : MUX2_X1 port map( A => n94, B => n83, S => A(23), Z => n65);
   U104 : NAND3_X1 port map( A1 => n66, A2 => n90, A3 => n65, ZN => p(23));
   U105 : MUX2_X1 port map( A => n80, B => n16, S => A(23), Z => n68);
   U106 : MUX2_X1 port map( A => n94, B => n83, S => n99, Z => n67);
   U107 : NAND3_X1 port map( A1 => n68, A2 => n90, A3 => n67, ZN => p(24));
   U108 : MUX2_X1 port map( A => n94, B => n83, S => n99, Z => n70);
   U109 : MUX2_X1 port map( A => n80, B => n16, S => n99, Z => n69);
   U110 : NAND3_X1 port map( A1 => n90, A2 => n70, A3 => n69, ZN => p(25));
   U111 : MUX2_X1 port map( A => n98, B => n16, S => n99, Z => n77);
   U112 : NAND3_X1 port map( A1 => n77, A2 => n76, A3 => n90, ZN => p(26));
   U113 : MUX2_X1 port map( A => n80, B => n16, S => n99, Z => n79);
   U114 : MUX2_X1 port map( A => n94, B => n83, S => n99, Z => n78);
   U115 : NAND3_X1 port map( A1 => n79, A2 => n90, A3 => n78, ZN => p(27));
   U116 : MUX2_X1 port map( A => n80, B => n16, S => n99, Z => n82);
   U117 : MUX2_X1 port map( A => n94, B => n83, S => n99, Z => n81);
   U118 : NAND3_X1 port map( A1 => n82, A2 => n90, A3 => n81, ZN => p(28));
   U119 : MUX2_X1 port map( A => n98, B => n16, S => n99, Z => n85);
   U120 : MUX2_X1 port map( A => n94, B => n83, S => n99, Z => n84);
   U121 : NAND3_X1 port map( A1 => n85, A2 => n90, A3 => n84, ZN => p(29));
   U122 : MUX2_X1 port map( A => n98, B => n16, S => n99, Z => n87);
   U123 : MUX2_X1 port map( A => n94, B => n88, S => n99, Z => n86);
   U124 : NAND3_X1 port map( A1 => n87, A2 => n90, A3 => n86, ZN => p(30));
   U125 : MUX2_X1 port map( A => n98, B => n16, S => n99, Z => n91);
   U126 : MUX2_X1 port map( A => n94, B => n4, S => n99, Z => n89);
   U127 : NAND3_X1 port map( A1 => n91, A2 => n90, A3 => n89, ZN => p(31));
   U128 : MUX2_X1 port map( A => n98, B => n16, S => n99, Z => n93);
   U129 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => p(32));
   U26 : INV_X1 port map( A => b(1), ZN => n47);
   U23 : INV_X1 port map( A => b(2), ZN => n71);
   U3 : NAND2_X1 port map( A1 => n96, A2 => n71, ZN => n4);
   U34 : NAND2_X2 port map( A1 => n17, A2 => b(2), ZN => n90);
   U35 : NAND2_X2 port map( A1 => b(2), A2 => n74, ZN => n94);
   U6 : INV_X1 port map( A => n72, ZN => n96);
   U7 : NAND3_X1 port map( A1 => n18, A2 => n47, A3 => b(2), ZN => n98);
   n99 <= '0';
   U5 : NAND2_X2 port map( A1 => b(1), A2 => b(0), ZN => n16);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_16 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_16;

architecture SYN_beh of ENC_16 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net32765, net32771, net32773, net32785, net32838, net32840, net32841,
      net33864, net33917, net32839, net32769, net32768, net32767, net32766, 
      net32786, net32794, net32764, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n69, n70, n71 : std_logic;

begin
   
   U6 : MUX2_X1 port map( A => net32764, B => net32771, S => n71, Z => n1);
   U7 : NAND3_X1 port map( A1 => net32768, A2 => net32769, A3 => n1, ZN => 
                           p(31));
   U9 : NAND2_X1 port map( A1 => n70, A2 => net32794, ZN => net32771);
   U10 : INV_X1 port map( A => b(2), ZN => net32794);
   U11 : NAND2_X1 port map( A1 => net32794, A2 => net33917, ZN => net33864);
   U12 : MUX2_X1 port map( A => net32794, B => n69, S => A(0), Z => n2);
   U13 : OAI211_X1 port map( C1 => net32794, C2 => net32841, A => net32766, B 
                           => n2, ZN => p(0));
   U14 : MUX2_X1 port map( A => net32766, B => net32767, S => n71, Z => 
                           net32765);
   U19 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => net32841);
   U23 : INV_X1 port map( A => b(0), ZN => net32839);
   U24 : XNOR2_X1 port map( A => b(0), B => net32838, ZN => net33917);
   U26 : MUX2_X1 port map( A => net32766, B => net32767, S => n71, Z => 
                           net32768);
   U32 : MUX2_X1 port map( A => net32764, B => net32771, S => n71, Z => 
                           net32773);
   U39 : MUX2_X1 port map( A => net32766, B => net32767, S => A(0), Z => n6);
   U40 : INV_X1 port map( A => net32841, ZN => net32840);
   U41 : MUX2_X1 port map( A => net32764, B => net33864, S => A(1), Z => n5);
   U42 : NAND3_X1 port map( A1 => n6, A2 => n4, A3 => n5, ZN => p(1));
   U43 : MUX2_X1 port map( A => net32766, B => net32767, S => A(1), Z => n8);
   U44 : MUX2_X1 port map( A => net32764, B => n69, S => A(2), Z => n7);
   U45 : NAND3_X1 port map( A1 => n8, A2 => net32769, A3 => n7, ZN => p(2));
   U46 : MUX2_X1 port map( A => net32766, B => net32767, S => A(2), Z => n10);
   U47 : MUX2_X1 port map( A => net32764, B => net33864, S => A(3), Z => n9);
   U48 : NAND3_X1 port map( A1 => n10, A2 => net32769, A3 => n9, ZN => p(3));
   U49 : MUX2_X1 port map( A => net32766, B => net32767, S => A(3), Z => n12);
   U50 : MUX2_X1 port map( A => net32764, B => n69, S => A(4), Z => n11);
   U51 : NAND3_X1 port map( A1 => n12, A2 => net32769, A3 => n11, ZN => p(4));
   U52 : MUX2_X1 port map( A => net32766, B => net32767, S => A(4), Z => n14);
   U53 : MUX2_X1 port map( A => net32764, B => net33864, S => A(5), Z => n13);
   U54 : NAND3_X1 port map( A1 => n14, A2 => net32769, A3 => n13, ZN => p(5));
   U55 : MUX2_X1 port map( A => net32766, B => net32767, S => A(5), Z => n16);
   U56 : MUX2_X1 port map( A => net32764, B => n69, S => A(6), Z => n15);
   U57 : NAND3_X1 port map( A1 => n16, A2 => net32769, A3 => n15, ZN => p(6));
   U58 : MUX2_X1 port map( A => net32766, B => net32767, S => A(6), Z => n18);
   U59 : MUX2_X1 port map( A => net32764, B => n69, S => A(7), Z => n17);
   U60 : NAND3_X1 port map( A1 => n18, A2 => net32769, A3 => n17, ZN => p(7));
   U61 : MUX2_X1 port map( A => net32766, B => net32767, S => A(7), Z => n20);
   U62 : MUX2_X1 port map( A => net32764, B => n69, S => A(8), Z => n19);
   U63 : NAND3_X1 port map( A1 => n19, A2 => net32769, A3 => n20, ZN => p(8));
   U64 : MUX2_X1 port map( A => net32766, B => net32767, S => A(8), Z => n22);
   U65 : MUX2_X1 port map( A => net32764, B => net33864, S => A(9), Z => n21);
   U66 : NAND3_X1 port map( A1 => n22, A2 => net32769, A3 => n21, ZN => p(9));
   U67 : MUX2_X1 port map( A => net32766, B => net32767, S => A(9), Z => n24);
   U68 : MUX2_X1 port map( A => net32764, B => n69, S => A(10), Z => n23);
   U69 : NAND3_X1 port map( A1 => n23, A2 => net32769, A3 => n24, ZN => p(10));
   U70 : MUX2_X1 port map( A => net32764, B => net33864, S => A(11), Z => n26);
   U71 : MUX2_X1 port map( A => net32766, B => net32767, S => A(10), Z => n25);
   U72 : NAND3_X1 port map( A1 => n26, A2 => net32769, A3 => n25, ZN => p(11));
   U73 : MUX2_X1 port map( A => net32766, B => net32767, S => A(11), Z => n28);
   U74 : MUX2_X1 port map( A => net32764, B => n69, S => A(12), Z => n27);
   U75 : NAND3_X1 port map( A1 => n28, A2 => net32769, A3 => n27, ZN => p(12));
   U76 : MUX2_X1 port map( A => net32764, B => net33864, S => A(13), Z => n30);
   U77 : MUX2_X1 port map( A => net32766, B => net32767, S => A(12), Z => n29);
   U78 : NAND3_X1 port map( A1 => net32769, A2 => n30, A3 => n29, ZN => p(13));
   U79 : MUX2_X1 port map( A => net32766, B => net32767, S => A(13), Z => n32);
   U80 : MUX2_X1 port map( A => net32764, B => net33864, S => A(14), Z => n31);
   U81 : NAND3_X1 port map( A1 => n32, A2 => net32769, A3 => n31, ZN => p(14));
   U82 : MUX2_X1 port map( A => net32766, B => net32767, S => A(14), Z => n34);
   U83 : MUX2_X1 port map( A => net32764, B => net33864, S => A(15), Z => n33);
   U84 : NAND3_X1 port map( A1 => n34, A2 => net32769, A3 => n33, ZN => p(15));
   U85 : MUX2_X1 port map( A => net32766, B => net32767, S => A(15), Z => n36);
   U86 : MUX2_X1 port map( A => net32764, B => n69, S => A(16), Z => n35);
   U87 : NAND3_X1 port map( A1 => n36, A2 => net32769, A3 => n35, ZN => p(16));
   U88 : MUX2_X1 port map( A => net32766, B => net32767, S => A(16), Z => n38);
   U89 : MUX2_X1 port map( A => net32764, B => net33864, S => A(17), Z => n37);
   U90 : NAND3_X1 port map( A1 => n38, A2 => net32769, A3 => n37, ZN => p(17));
   U91 : MUX2_X1 port map( A => net32766, B => net32767, S => A(17), Z => n40);
   U92 : MUX2_X1 port map( A => net32764, B => n69, S => A(18), Z => n39);
   U93 : NAND3_X1 port map( A1 => n40, A2 => net32769, A3 => n39, ZN => p(18));
   U94 : MUX2_X1 port map( A => net32766, B => net32767, S => A(18), Z => n42);
   U95 : MUX2_X1 port map( A => net32764, B => n69, S => A(19), Z => n41);
   U96 : NAND3_X1 port map( A1 => n42, A2 => net32769, A3 => n41, ZN => p(19));
   U97 : MUX2_X1 port map( A => net32766, B => net32767, S => A(19), Z => n44);
   U98 : MUX2_X1 port map( A => net32764, B => net33864, S => A(20), Z => n43);
   U99 : NAND3_X1 port map( A1 => n44, A2 => n4, A3 => n43, ZN => p(20));
   U100 : MUX2_X1 port map( A => net32766, B => net32767, S => A(20), Z => n46)
                           ;
   U101 : MUX2_X1 port map( A => net32764, B => net33864, S => A(21), Z => n45)
                           ;
   U102 : NAND3_X1 port map( A1 => n46, A2 => n4, A3 => n45, ZN => p(21));
   U103 : MUX2_X1 port map( A => net32766, B => net32767, S => A(21), Z => n48)
                           ;
   U104 : MUX2_X1 port map( A => net32764, B => net32771, S => A(22), Z => n47)
                           ;
   U105 : NAND3_X1 port map( A1 => n48, A2 => n4, A3 => n47, ZN => p(22));
   U106 : MUX2_X1 port map( A => net32766, B => net32767, S => A(22), Z => n50)
                           ;
   U107 : MUX2_X1 port map( A => net32764, B => net32771, S => A(23), Z => n49)
                           ;
   U108 : NAND3_X1 port map( A1 => n50, A2 => n4, A3 => n49, ZN => p(23));
   U109 : MUX2_X1 port map( A => net32766, B => net32767, S => A(23), Z => n52)
                           ;
   U110 : MUX2_X1 port map( A => net32764, B => net32771, S => n71, Z => n51);
   U111 : NAND3_X1 port map( A1 => n52, A2 => n4, A3 => n51, ZN => p(24));
   U112 : MUX2_X1 port map( A => net32766, B => net32767, S => n71, Z => n55);
   U113 : INV_X1 port map( A => net32786, ZN => net32785);
   U116 : NAND3_X1 port map( A1 => n54, A2 => n4, A3 => n55, ZN => p(25));
   U117 : MUX2_X1 port map( A => net32766, B => net32767, S => n71, Z => n57);
   U118 : MUX2_X1 port map( A => net32764, B => net32771, S => n71, Z => n56);
   U119 : NAND3_X1 port map( A1 => n56, A2 => n4, A3 => n57, ZN => p(26));
   U120 : MUX2_X1 port map( A => net32766, B => net32841, S => n71, Z => n59);
   U121 : MUX2_X1 port map( A => net32764, B => net32771, S => n71, Z => n58);
   U122 : NAND3_X1 port map( A1 => n58, A2 => n4, A3 => n59, ZN => p(27));
   U123 : MUX2_X1 port map( A => net32766, B => net32767, S => n71, Z => n61);
   U124 : MUX2_X1 port map( A => net32764, B => net32771, S => n71, Z => n60);
   U125 : NAND3_X1 port map( A1 => n61, A2 => n4, A3 => n60, ZN => p(28));
   U126 : MUX2_X1 port map( A => net32766, B => net32767, S => n71, Z => n63);
   U127 : MUX2_X1 port map( A => net32764, B => net32771, S => n71, Z => n62);
   U128 : NAND3_X1 port map( A1 => n63, A2 => n4, A3 => n62, ZN => p(29));
   U129 : MUX2_X1 port map( A => net32766, B => net32767, S => n71, Z => n64);
   U130 : NAND3_X1 port map( A1 => n64, A2 => n4, A3 => net32773, ZN => p(30));
   U131 : NAND2_X1 port map( A1 => net32765, A2 => net32764, ZN => p(32));
   U20 : INV_X1 port map( A => b(1), ZN => net32838);
   U18 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => net32786);
   U15 : NAND2_X2 port map( A1 => b(2), A2 => net32786, ZN => net32764);
   U29 : NAND2_X1 port map( A1 => net32840, A2 => b(2), ZN => net32769);
   U8 : NAND2_X1 port map( A1 => net32840, A2 => b(2), ZN => n4);
   U16 : NAND2_X1 port map( A1 => net32785, A2 => net32771, ZN => n53);
   U17 : NAND2_X1 port map( A1 => net32794, A2 => n70, ZN => n69);
   U22 : NAND2_X1 port map( A1 => b(2), A2 => n53, ZN => n54);
   U25 : XNOR2_X1 port map( A => b(0), B => net32838, ZN => n70);
   n71 <= '0';
   U3 : NAND3_X2 port map( A1 => b(2), A2 => net32839, A3 => net32838, ZN => 
                           net32766);
   U4 : NAND2_X2 port map( A1 => b(0), A2 => b(1), ZN => net32767);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_0 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_0;

architecture SYN_beh of ENC_0 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n72, n73, n75, n77, n79, n81
      , n82, n86, n88, n93, n96, n97, n98, n99, n100, n101, n102, n103, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n118, 
      n120, n121, n122, n123, n124 : std_logic;

begin
   
   U19 : INV_X1 port map( A => b(2), ZN => n19);
   U25 : MUX2_X1 port map( A => n19, B => n81, S => A(0), Z => n18);
   U26 : OAI211_X1 port map( C1 => n19, C2 => n123, A => n86, B => n18, ZN => 
                           p(0));
   U30 : MUX2_X1 port map( A => n88, B => n81, S => A(1), Z => n21);
   U33 : MUX2_X1 port map( A => n88, B => n81, S => A(2), Z => n23);
   U36 : MUX2_X1 port map( A => n88, B => n81, S => A(3), Z => n25);
   U39 : MUX2_X1 port map( A => n88, B => n81, S => A(4), Z => n27);
   U42 : MUX2_X1 port map( A => n88, B => n81, S => A(5), Z => n29);
   U45 : MUX2_X1 port map( A => n88, B => n81, S => A(6), Z => n31);
   U48 : MUX2_X1 port map( A => n88, B => n81, S => A(7), Z => n33);
   U51 : MUX2_X1 port map( A => n88, B => n81, S => A(8), Z => n35);
   U54 : MUX2_X1 port map( A => n88, B => n81, S => A(9), Z => n37);
   U57 : MUX2_X1 port map( A => n88, B => n81, S => A(10), Z => n39);
   U60 : MUX2_X1 port map( A => n88, B => n81, S => A(11), Z => n41);
   U63 : MUX2_X1 port map( A => n88, B => n81, S => A(12), Z => n43);
   U66 : MUX2_X1 port map( A => n88, B => n81, S => A(13), Z => n45);
   U69 : MUX2_X1 port map( A => n88, B => n81, S => A(14), Z => n47);
   U71 : MUX2_X1 port map( A => n88, B => n81, S => A(15), Z => n50);
   U75 : MUX2_X1 port map( A => n88, B => n81, S => A(16), Z => n51);
   U78 : MUX2_X1 port map( A => n88, B => n81, S => A(17), Z => n53);
   U81 : MUX2_X1 port map( A => n88, B => n81, S => A(18), Z => n55);
   U84 : MUX2_X1 port map( A => n88, B => n81, S => A(19), Z => n57);
   U87 : MUX2_X1 port map( A => n88, B => n81, S => A(20), Z => n59);
   U90 : MUX2_X1 port map( A => n88, B => n81, S => A(21), Z => n61);
   U93 : MUX2_X1 port map( A => n88, B => n81, S => A(22), Z => n63);
   U95 : MUX2_X1 port map( A => n88, B => n81, S => A(23), Z => n66);
   U99 : MUX2_X1 port map( A => n88, B => n81, S => n124, Z => n67);
   U102 : MUX2_X1 port map( A => n88, B => n81, S => n124, Z => n69);
   U104 : MUX2_X1 port map( A => n88, B => n81, S => n124, Z => n72);
   U108 : MUX2_X1 port map( A => n88, B => n81, S => n124, Z => n73);
   U111 : MUX2_X1 port map( A => n88, B => n81, S => n124, Z => n75);
   U114 : MUX2_X1 port map( A => n88, B => n81, S => n124, Z => n77);
   U117 : MUX2_X1 port map( A => n88, B => n81, S => n124, Z => n79);
   U120 : MUX2_X1 port map( A => n88, B => n81, S => n124, Z => n82);
   U123 : NAND2_X1 port map( A1 => n88, A2 => n86, ZN => p(32));
   U5 : NAND2_X1 port map( A1 => n86, A2 => n82, ZN => p(31));
   U7 : NAND2_X1 port map( A1 => n48, A2 => n47, ZN => p(14));
   U8 : NAND2_X1 port map( A1 => n46, A2 => n45, ZN => p(13));
   U9 : NAND2_X1 port map( A1 => n36, A2 => n35, ZN => p(8));
   U10 : NAND2_X1 port map( A1 => n32, A2 => n31, ZN => p(6));
   U11 : NAND2_X1 port map( A1 => n28, A2 => n27, ZN => p(4));
   U12 : NAND2_X1 port map( A1 => n93, A2 => n113, ZN => n62);
   U13 : NAND2_X1 port map( A1 => n93, A2 => n110, ZN => n68);
   U14 : NAND2_X1 port map( A1 => n93, A2 => n107, ZN => n26);
   U15 : INV_X1 port map( A => A(19), ZN => n114);
   U16 : INV_X1 port map( A => A(16), ZN => n118);
   U17 : INV_X1 port map( A => A(15), ZN => n120);
   U20 : INV_X1 port map( A => A(2), ZN => n107);
   U21 : INV_X1 port map( A => A(21), ZN => n112);
   U22 : NAND2_X1 port map( A1 => b(1), A2 => b(2), ZN => n88);
   U23 : INV_X1 port map( A => A(20), ZN => n113);
   U24 : INV_X1 port map( A => A(17), ZN => n116);
   U27 : INV_X1 port map( A => A(22), ZN => n111);
   U28 : NAND2_X1 port map( A1 => n93, A2 => n108, ZN => n24);
   U29 : NAND2_X1 port map( A1 => n93, A2 => n122, ZN => n48);
   U31 : NAND2_X1 port map( A1 => n93, A2 => n111, ZN => n65);
   U32 : NAND2_X1 port map( A1 => n93, A2 => n112, ZN => n64);
   U34 : INV_X1 port map( A => A(18), ZN => n115);
   U35 : NAND2_X1 port map( A1 => n24, A2 => n23, ZN => p(2));
   U37 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => p(22));
   U38 : NAND2_X1 port map( A1 => n93, A2 => n121, ZN => n49);
   U40 : NAND2_X1 port map( A1 => n93, A2 => n97, ZN => n44);
   U41 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => p(21));
   U43 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => p(15));
   U44 : NAND2_X1 port map( A1 => n44, A2 => n43, ZN => p(12));
   U46 : NAND2_X1 port map( A1 => n68, A2 => n67, ZN => p(24));
   U47 : NAND2_X1 port map( A1 => n58, A2 => n57, ZN => p(19));
   U49 : NAND2_X1 port map( A1 => n52, A2 => n51, ZN => p(16));
   U50 : NAND2_X1 port map( A1 => n56, A2 => n55, ZN => p(18));
   U52 : NAND2_X1 port map( A1 => n26, A2 => n25, ZN => p(3));
   U53 : NAND2_X1 port map( A1 => n30, A2 => n29, ZN => p(5));
   U55 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => p(7));
   U56 : NAND2_X1 port map( A1 => n60, A2 => n59, ZN => p(20));
   U59 : INV_X1 port map( A => b(1), ZN => n17);
   U61 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => p(23));
   U62 : INV_X1 port map( A => A(23), ZN => n110);
   U64 : NAND2_X1 port map( A1 => n72, A2 => n86, ZN => p(26));
   U65 : NAND2_X1 port map( A1 => n86, A2 => n79, ZN => p(30));
   U67 : NAND2_X1 port map( A1 => n86, A2 => n77, ZN => p(29));
   U68 : NAND2_X1 port map( A1 => n86, A2 => n69, ZN => p(25));
   U70 : NAND2_X1 port map( A1 => n86, A2 => n73, ZN => p(27));
   U72 : NAND2_X1 port map( A1 => n86, A2 => n75, ZN => p(28));
   U76 : NAND2_X1 port map( A1 => n22, A2 => n21, ZN => p(1));
   U77 : NAND2_X1 port map( A1 => n54, A2 => n53, ZN => p(17));
   U79 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => p(11));
   U80 : NAND2_X1 port map( A1 => n40, A2 => n39, ZN => p(10));
   U82 : NAND2_X1 port map( A1 => n38, A2 => n37, ZN => p(9));
   U83 : NAND2_X1 port map( A1 => n93, A2 => n96, ZN => n46);
   U85 : INV_X1 port map( A => A(12), ZN => n96);
   U86 : INV_X1 port map( A => A(11), ZN => n97);
   U88 : NAND2_X1 port map( A1 => n93, A2 => n98, ZN => n42);
   U89 : INV_X1 port map( A => A(10), ZN => n98);
   U91 : NAND2_X1 port map( A1 => n93, A2 => n99, ZN => n40);
   U92 : INV_X1 port map( A => A(9), ZN => n99);
   U94 : NAND2_X1 port map( A1 => n93, A2 => n100, ZN => n38);
   U96 : INV_X1 port map( A => A(8), ZN => n100);
   U97 : NAND2_X1 port map( A1 => n93, A2 => n101, ZN => n36);
   U98 : INV_X1 port map( A => A(7), ZN => n101);
   U100 : NAND2_X1 port map( A1 => n93, A2 => n102, ZN => n34);
   U101 : INV_X1 port map( A => A(6), ZN => n102);
   U103 : NAND2_X1 port map( A1 => n93, A2 => n103, ZN => n32);
   U105 : INV_X1 port map( A => A(5), ZN => n103);
   U106 : NAND2_X1 port map( A1 => n93, A2 => n105, ZN => n30);
   U107 : INV_X1 port map( A => A(4), ZN => n105);
   U109 : NAND2_X1 port map( A1 => n93, A2 => n106, ZN => n28);
   U110 : INV_X1 port map( A => A(3), ZN => n106);
   U112 : INV_X1 port map( A => A(1), ZN => n108);
   U113 : NAND2_X1 port map( A1 => n93, A2 => n109, ZN => n22);
   U115 : INV_X1 port map( A => A(0), ZN => n109);
   U116 : NAND2_X1 port map( A1 => n93, A2 => n114, ZN => n60);
   U118 : NAND2_X1 port map( A1 => n93, A2 => n115, ZN => n58);
   U119 : NAND2_X1 port map( A1 => n93, A2 => n116, ZN => n56);
   U121 : NAND2_X1 port map( A1 => n93, A2 => n118, ZN => n54);
   U122 : NAND2_X1 port map( A1 => n93, A2 => n120, ZN => n52);
   U124 : INV_X1 port map( A => A(14), ZN => n121);
   U125 : INV_X1 port map( A => A(13), ZN => n122);
   n123 <= '1';
   n124 <= '0';
   U3 : OR2_X2 port map( A1 => b(2), A2 => n17, ZN => n81);
   U4 : NAND2_X2 port map( A1 => n17, A2 => b(2), ZN => n86);
   U6 : INV_X2 port map( A => n86, ZN => n93);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PackFP is

   port( SIGN : in std_logic;  EXP : in std_logic_vector (7 downto 0);  SIG : 
         in std_logic_vector (22 downto 0);  isNaN, isINF, isZ : in std_logic; 
         FP : out std_logic_vector (31 downto 0);  clk : in std_logic);

end PackFP;

architecture SYN_PackFP of PackFP is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal FP_30_port, FP_29_port, FP_28_port, FP_27_port, FP_26_port, 
      FP_25_port, FP_24_port, FP_23_port, FP_22_port, FP_21_port, FP_20_port, 
      FP_19_port, FP_18_port, FP_17_port, FP_16_port, FP_15_port, FP_14_port, 
      FP_13_port, FP_12_port, FP_11_port, FP_10_port, FP_9_port, FP_8_port, 
      FP_7_port, FP_6_port, FP_5_port, FP_4_port, FP_3_port, FP_2_port, 
      FP_1_port, FP_0_port, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n18, n19, n21, n22, n23, n_2133 : std_logic;

begin
   FP <= ( SIGN, FP_30_port, FP_29_port, FP_28_port, FP_27_port, FP_26_port, 
      FP_25_port, FP_24_port, FP_23_port, FP_22_port, FP_21_port, FP_20_port, 
      FP_19_port, FP_18_port, FP_17_port, FP_16_port, FP_15_port, FP_14_port, 
      FP_13_port, FP_12_port, FP_11_port, FP_10_port, FP_9_port, FP_8_port, 
      FP_7_port, FP_6_port, FP_5_port, FP_4_port, FP_3_port, FP_2_port, 
      FP_1_port, FP_0_port );
   
   U7 : INV_X1 port map( A => isNaN, ZN => n5);
   U9 : AND2_X1 port map( A1 => SIG(0), A2 => n23, ZN => FP_0_port);
   U10 : AND2_X1 port map( A1 => SIG(1), A2 => n23, ZN => FP_1_port);
   U11 : AND2_X1 port map( A1 => SIG(2), A2 => n23, ZN => FP_2_port);
   U12 : AND2_X1 port map( A1 => SIG(3), A2 => n23, ZN => FP_3_port);
   U13 : AND2_X1 port map( A1 => SIG(4), A2 => n23, ZN => FP_4_port);
   U14 : AND2_X1 port map( A1 => SIG(5), A2 => n23, ZN => FP_5_port);
   U15 : AND2_X1 port map( A1 => SIG(6), A2 => n23, ZN => FP_6_port);
   U16 : AND2_X1 port map( A1 => n23, A2 => SIG(7), ZN => FP_7_port);
   U17 : AND2_X1 port map( A1 => n23, A2 => SIG(8), ZN => FP_8_port);
   U18 : AND2_X1 port map( A1 => SIG(9), A2 => n23, ZN => FP_9_port);
   U19 : AND2_X1 port map( A1 => SIG(10), A2 => n23, ZN => FP_10_port);
   U20 : AND2_X1 port map( A1 => SIG(11), A2 => n1, ZN => FP_11_port);
   U21 : AND2_X1 port map( A1 => n1, A2 => SIG(12), ZN => FP_12_port);
   U22 : AND2_X1 port map( A1 => n1, A2 => SIG(13), ZN => FP_13_port);
   U23 : AND2_X1 port map( A1 => n1, A2 => SIG(14), ZN => FP_14_port);
   U24 : AND2_X1 port map( A1 => SIG(15), A2 => n1, ZN => FP_15_port);
   U25 : AND2_X1 port map( A1 => SIG(16), A2 => n1, ZN => FP_16_port);
   U26 : AND2_X1 port map( A1 => SIG(17), A2 => n1, ZN => FP_17_port);
   U27 : AND2_X1 port map( A1 => SIG(18), A2 => n1, ZN => FP_18_port);
   U28 : AND2_X1 port map( A1 => SIG(19), A2 => n1, ZN => FP_19_port);
   U29 : AND2_X1 port map( A1 => SIG(20), A2 => n1, ZN => FP_20_port);
   U30 : AND2_X1 port map( A1 => n1, A2 => SIG(21), ZN => FP_21_port);
   U31 : NAND3_X1 port map( A1 => n3, A2 => SIG(22), A3 => n14, ZN => n4);
   U32 : NAND2_X1 port map( A1 => n4, A2 => n18, ZN => FP_22_port);
   U33 : AOI21_X1 port map( B1 => EXP(0), B2 => n14, A => n13, ZN => n6);
   U34 : INV_X1 port map( A => n6, ZN => FP_23_port);
   U35 : AOI21_X1 port map( B1 => EXP(1), B2 => n14, A => n13, ZN => n7);
   U36 : INV_X1 port map( A => n7, ZN => FP_24_port);
   U37 : AOI21_X1 port map( B1 => EXP(2), B2 => n14, A => n13, ZN => n8);
   U38 : INV_X1 port map( A => n8, ZN => FP_25_port);
   U39 : AOI21_X1 port map( B1 => EXP(3), B2 => n14, A => n13, ZN => n9);
   U40 : INV_X1 port map( A => n9, ZN => FP_26_port);
   U41 : AOI21_X1 port map( B1 => EXP(4), B2 => n14, A => n13, ZN => n10);
   U42 : INV_X1 port map( A => n10, ZN => FP_27_port);
   U43 : AOI21_X1 port map( B1 => EXP(5), B2 => n14, A => n13, ZN => n11);
   U44 : INV_X1 port map( A => n11, ZN => FP_28_port);
   U45 : AOI21_X1 port map( B1 => EXP(6), B2 => n14, A => n13, ZN => n12);
   U46 : INV_X1 port map( A => n12, ZN => FP_29_port);
   U47 : AOI21_X1 port map( B1 => EXP(7), B2 => n14, A => n13, ZN => n15);
   U48 : INV_X1 port map( A => n15, ZN => FP_30_port);
   U5 : INV_X1 port map( A => isZ, ZN => n14);
   U3 : NOR2_X2 port map( A1 => isINF, A2 => n21, ZN => n22);
   U4 : OR2_X2 port map( A1 => isINF, A2 => n21, ZN => n13);
   U8 : INV_X1 port map( A => isINF, ZN => n3);
   U49 : AND2_X2 port map( A1 => n22, A2 => n14, ZN => n23);
   U50 : AND2_X2 port map( A1 => n22, A2 => n14, ZN => n1);
   MY_CLK_r_REG7_S4 : DFF_X1 port map( D => n19, CK => clk, Q => n18, QN => n21
                           );
   MY_CLK_r_REG6_S3 : DFF_X1 port map( D => n5, CK => clk, Q => n19, QN => 
                           n_2133);

end SYN_PackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPnormalize_SIG_width28_1 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
         std_logic);

end FPnormalize_SIG_width28_1;

architecture SYN_FPnormalize of FPnormalize_SIG_width28_1 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n6, n7, n8, n9, n10, n11, n13, n14, n16, n20, n28, n29, n30, n31,
      n32, n33, n34, n35, n37, n41, n42, n43, n44, n45, n46, n47, n_2141, 
      n_2142, n_2143, n_2144, n_2145, n_2146 : std_logic;

begin
   
   U4 : INV_X1 port map( A => SIG_in(27), ZN => n4);
   U9 : XOR2_X1 port map( A => n29, B => SIG_in(27), Z => EXP_out(0));
   U11 : NOR2_X1 port map( A1 => n4, A2 => n42, ZN => n6);
   U12 : XOR2_X1 port map( A => n30, B => n6, Z => EXP_out(1));
   U13 : NAND3_X1 port map( A1 => n30, A2 => SIG_in(27), A3 => n29, ZN => n7);
   U14 : INV_X1 port map( A => n7, ZN => n10);
   U15 : XOR2_X1 port map( A => n31, B => n37, Z => EXP_out(2));
   U16 : INV_X1 port map( A => EXP_in(2), ZN => n8);
   U17 : NOR2_X1 port map( A1 => n7, A2 => n8, ZN => n9);
   U18 : XOR2_X1 port map( A => n32, B => n28, Z => EXP_out(3));
   U19 : NAND3_X1 port map( A1 => n32, A2 => n31, A3 => n37, ZN => n11);
   U20 : INV_X1 port map( A => n11, ZN => n14);
   U23 : NOR2_X1 port map( A1 => n46, A2 => n11, ZN => n13);
   U33 : MUX2_X1 port map( A => SIG_in(3), B => SIG_in(4), S => SIG_in(27), Z 
                           => SIG_out(3));
   U34 : MUX2_X1 port map( A => SIG_in(4), B => SIG_in(5), S => SIG_in(27), Z 
                           => SIG_out(4));
   U35 : MUX2_X1 port map( A => SIG_in(5), B => SIG_in(6), S => SIG_in(27), Z 
                           => SIG_out(5));
   U36 : MUX2_X1 port map( A => SIG_in(6), B => SIG_in(7), S => SIG_in(27), Z 
                           => SIG_out(6));
   U37 : MUX2_X1 port map( A => SIG_in(7), B => SIG_in(8), S => SIG_in(27), Z 
                           => SIG_out(7));
   U38 : MUX2_X1 port map( A => SIG_in(8), B => SIG_in(9), S => SIG_in(27), Z 
                           => SIG_out(8));
   U39 : MUX2_X1 port map( A => SIG_in(9), B => SIG_in(10), S => SIG_in(27), Z 
                           => SIG_out(9));
   U40 : MUX2_X1 port map( A => SIG_in(10), B => SIG_in(11), S => SIG_in(27), Z
                           => SIG_out(10));
   U41 : MUX2_X1 port map( A => SIG_in(11), B => SIG_in(12), S => SIG_in(27), Z
                           => SIG_out(11));
   U42 : MUX2_X1 port map( A => SIG_in(12), B => SIG_in(13), S => SIG_in(27), Z
                           => SIG_out(12));
   U43 : MUX2_X1 port map( A => SIG_in(13), B => SIG_in(14), S => SIG_in(27), Z
                           => SIG_out(13));
   U44 : MUX2_X1 port map( A => SIG_in(14), B => SIG_in(15), S => SIG_in(27), Z
                           => SIG_out(14));
   U45 : MUX2_X1 port map( A => SIG_in(15), B => SIG_in(16), S => SIG_in(27), Z
                           => SIG_out(15));
   U46 : MUX2_X1 port map( A => SIG_in(16), B => SIG_in(17), S => SIG_in(27), Z
                           => SIG_out(16));
   U47 : MUX2_X1 port map( A => SIG_in(17), B => SIG_in(18), S => SIG_in(27), Z
                           => SIG_out(17));
   U48 : MUX2_X1 port map( A => SIG_in(18), B => SIG_in(19), S => SIG_in(27), Z
                           => SIG_out(18));
   U49 : MUX2_X1 port map( A => SIG_in(19), B => SIG_in(20), S => SIG_in(27), Z
                           => SIG_out(19));
   U50 : MUX2_X1 port map( A => SIG_in(20), B => SIG_in(21), S => SIG_in(27), Z
                           => SIG_out(20));
   U51 : MUX2_X1 port map( A => SIG_in(21), B => SIG_in(22), S => SIG_in(27), Z
                           => SIG_out(21));
   U52 : MUX2_X1 port map( A => SIG_in(22), B => SIG_in(23), S => SIG_in(27), Z
                           => SIG_out(22));
   U53 : MUX2_X1 port map( A => SIG_in(23), B => SIG_in(24), S => SIG_in(27), Z
                           => SIG_out(23));
   U54 : MUX2_X1 port map( A => SIG_in(24), B => SIG_in(25), S => SIG_in(27), Z
                           => SIG_out(24));
   U55 : MUX2_X1 port map( A => SIG_in(25), B => SIG_in(26), S => SIG_in(27), Z
                           => SIG_out(25));
   U56 : INV_X1 port map( A => SIG_in(26), ZN => n20);
   U57 : NAND2_X1 port map( A1 => n20, A2 => n4, ZN => SIG_out(26));
   MY_CLK_r_REG61_S4 : DFF_X1 port map( D => EXP_in(7), CK => clk, Q => n_2141,
                           QN => n43);
   U2 : OR2_X2 port map( A1 => n11, A2 => n47, ZN => n16);
   U3 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => n47);
   U5 : NOR2_X1 port map( A1 => n16, A2 => n44, ZN => n45);
   U6 : XNOR2_X1 port map( A => n45, B => n43, ZN => EXP_out(7));
   U7 : XNOR2_X1 port map( A => n14, B => n46, ZN => EXP_out(4));
   U8 : XNOR2_X1 port map( A => n16, B => n35, ZN => EXP_out(6));
   U10 : XNOR2_X1 port map( A => n13, B => n41, ZN => EXP_out(5));
   MY_CLK_r_REG66_S3 : DFF_X1 port map( D => EXP_in(0), CK => clk, Q => n29, QN
                           => n42);
   MY_CLK_r_REG63_S4 : DFF_X1 port map( D => EXP_in(4), CK => clk, Q => n33, QN
                           => n46);
   MY_CLK_r_REG62_S4 : DFF_X1 port map( D => EXP_in(6), CK => clk, Q => n35, QN
                           => n44);
   MY_CLK_r_REG60_S4 : DFF_X1 port map( D => EXP_in(5), CK => clk, Q => n34, QN
                           => n41);
   MY_CLK_r_REG65_S4 : DFF_X1 port map( D => EXP_in(3), CK => clk, Q => n32, QN
                           => n_2142);
   MY_CLK_r_REG64_S4 : DFF_X1 port map( D => EXP_in(2), CK => clk, Q => n31, QN
                           => n_2143);
   MY_CLK_r_REG21_S4 : DFF_X1 port map( D => n10, CK => clk, Q => n37, QN => 
                           n_2144);
   MY_CLK_r_REG20_S4 : DFF_X1 port map( D => n9, CK => clk, Q => n28, QN => 
                           n_2145);
   MY_CLK_r_REG18_S3 : DFF_X1 port map( D => EXP_in(1), CK => clk, Q => n30, QN
                           => n_2146);

end SYN_FPnormalize;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPround_SIG_width28 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
         std_logic);

end FPround_SIG_width28;

architecture SYN_FPround of FPround_SIG_width28 is

   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FPround_SIG_width28_DW01_inc_1
      port( A : in std_logic_vector (24 downto 0);  SUM : out std_logic_vector 
            (24 downto 0));
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n55, n58, n_2153, n_2154, n_2155, n_2156, n_2157
      , n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166,
      n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, 
      n_2176, n_2177 : std_logic;

begin
   EXP_out <= ( EXP_in(7), EXP_in(6), EXP_in(5), EXP_in(4), EXP_in(3), 
      EXP_in(2), EXP_in(1), EXP_in(0) );
   
   U8 : MUX2_X1 port map( A => n30, B => N2, S => n55, Z => SIG_out(3));
   U9 : MUX2_X1 port map( A => n31, B => N3, S => n55, Z => SIG_out(4));
   U10 : MUX2_X1 port map( A => n32, B => N4, S => n55, Z => SIG_out(5));
   U11 : MUX2_X1 port map( A => n33, B => N5, S => n55, Z => SIG_out(6));
   U12 : MUX2_X1 port map( A => n34, B => N6, S => n55, Z => SIG_out(7));
   U13 : MUX2_X1 port map( A => n35, B => N7, S => n55, Z => SIG_out(8));
   U14 : MUX2_X1 port map( A => n36, B => N8, S => n55, Z => SIG_out(9));
   U15 : MUX2_X1 port map( A => n37, B => N9, S => n55, Z => SIG_out(10));
   U16 : MUX2_X1 port map( A => n38, B => N10, S => n55, Z => SIG_out(11));
   U17 : MUX2_X1 port map( A => n39, B => N11, S => n55, Z => SIG_out(12));
   U18 : MUX2_X1 port map( A => n40, B => N12, S => n55, Z => SIG_out(13));
   U19 : MUX2_X1 port map( A => n41, B => N13, S => n55, Z => SIG_out(14));
   U20 : MUX2_X1 port map( A => n42, B => N14, S => n55, Z => SIG_out(15));
   U21 : MUX2_X1 port map( A => n43, B => N15, S => n55, Z => SIG_out(16));
   U22 : MUX2_X1 port map( A => n44, B => N16, S => n55, Z => SIG_out(17));
   U23 : MUX2_X1 port map( A => n45, B => N17, S => n55, Z => SIG_out(18));
   U24 : MUX2_X1 port map( A => n46, B => N18, S => n55, Z => SIG_out(19));
   U25 : MUX2_X1 port map( A => n47, B => N19, S => n55, Z => SIG_out(20));
   U26 : MUX2_X1 port map( A => n48, B => N20, S => n55, Z => SIG_out(21));
   U27 : MUX2_X1 port map( A => n49, B => N21, S => n55, Z => SIG_out(22));
   U28 : MUX2_X1 port map( A => n50, B => N22, S => n55, Z => SIG_out(23));
   U29 : MUX2_X1 port map( A => n51, B => N23, S => n55, Z => SIG_out(24));
   U30 : MUX2_X1 port map( A => n52, B => N24, S => n55, Z => SIG_out(25));
   U31 : MUX2_X1 port map( A => n53, B => N25, S => n55, Z => SIG_out(26));
   U4 : AND2_X2 port map( A1 => n55, A2 => N26, ZN => SIG_out(27));
   n58 <= '0';
   add_45 : FPround_SIG_width28_DW01_inc_1 port map( A(24) => n58, A(23) => n53
                           , A(22) => n52, A(21) => n51, A(20) => n50, A(19) =>
                           n49, A(18) => n48, A(17) => n47, A(16) => n46, A(15)
                           => n45, A(14) => n44, A(13) => n43, A(12) => n42, 
                           A(11) => n41, A(10) => n40, A(9) => n39, A(8) => n38
                           , A(7) => n37, A(6) => n36, A(5) => n35, A(4) => n34
                           , A(3) => n33, A(2) => n32, A(1) => n31, A(0) => n30
                           , SUM(24) => N26, SUM(23) => N25, SUM(22) => N24, 
                           SUM(21) => N23, SUM(20) => N22, SUM(19) => N21, 
                           SUM(18) => N20, SUM(17) => N19, SUM(16) => N18, 
                           SUM(15) => N17, SUM(14) => N16, SUM(13) => N15, 
                           SUM(12) => N14, SUM(11) => N13, SUM(10) => N12, 
                           SUM(9) => N11, SUM(8) => N10, SUM(7) => N9, SUM(6) 
                           => N8, SUM(5) => N7, SUM(4) => N6, SUM(3) => N5, 
                           SUM(2) => N4, SUM(1) => N3, SUM(0) => N2);
   MY_CLK_r_REG79_S3 : DFF_X1 port map( D => SIG_in(25), CK => clk, Q => n52, 
                           QN => n_2153);
   MY_CLK_r_REG78_S3 : DFF_X1 port map( D => SIG_in(13), CK => clk, Q => n40, 
                           QN => n_2154);
   MY_CLK_r_REG77_S3 : DFF_X1 port map( D => SIG_in(14), CK => clk, Q => n41, 
                           QN => n_2155);
   MY_CLK_r_REG76_S3 : DFF_X1 port map( D => SIG_in(15), CK => clk, Q => n42, 
                           QN => n_2156);
   MY_CLK_r_REG75_S3 : DFF_X1 port map( D => SIG_in(16), CK => clk, Q => n43, 
                           QN => n_2157);
   MY_CLK_r_REG74_S3 : DFF_X1 port map( D => SIG_in(17), CK => clk, Q => n44, 
                           QN => n_2158);
   MY_CLK_r_REG73_S3 : DFF_X1 port map( D => SIG_in(18), CK => clk, Q => n45, 
                           QN => n_2159);
   MY_CLK_r_REG72_S3 : DFF_X1 port map( D => SIG_in(19), CK => clk, Q => n46, 
                           QN => n_2160);
   MY_CLK_r_REG71_S3 : DFF_X1 port map( D => SIG_in(20), CK => clk, Q => n47, 
                           QN => n_2161);
   MY_CLK_r_REG70_S3 : DFF_X1 port map( D => SIG_in(21), CK => clk, Q => n48, 
                           QN => n_2162);
   MY_CLK_r_REG69_S3 : DFF_X1 port map( D => SIG_in(22), CK => clk, Q => n49, 
                           QN => n_2163);
   MY_CLK_r_REG68_S3 : DFF_X1 port map( D => SIG_in(23), CK => clk, Q => n50, 
                           QN => n_2164);
   MY_CLK_r_REG67_S3 : DFF_X1 port map( D => SIG_in(24), CK => clk, Q => n51, 
                           QN => n_2165);
   MY_CLK_r_REG57_S3 : DFF_X1 port map( D => SIG_in(3), CK => clk, Q => n30, QN
                           => n_2166);
   MY_CLK_r_REG56_S3 : DFF_X1 port map( D => SIG_in(4), CK => clk, Q => n31, QN
                           => n_2167);
   MY_CLK_r_REG55_S3 : DFF_X1 port map( D => SIG_in(5), CK => clk, Q => n32, QN
                           => n_2168);
   MY_CLK_r_REG54_S3 : DFF_X1 port map( D => SIG_in(6), CK => clk, Q => n33, QN
                           => n_2169);
   MY_CLK_r_REG53_S3 : DFF_X1 port map( D => SIG_in(7), CK => clk, Q => n34, QN
                           => n_2170);
   MY_CLK_r_REG52_S3 : DFF_X1 port map( D => SIG_in(8), CK => clk, Q => n35, QN
                           => n_2171);
   MY_CLK_r_REG51_S3 : DFF_X1 port map( D => SIG_in(9), CK => clk, Q => n36, QN
                           => n_2172);
   MY_CLK_r_REG50_S3 : DFF_X1 port map( D => SIG_in(10), CK => clk, Q => n37, 
                           QN => n_2173);
   MY_CLK_r_REG49_S3 : DFF_X1 port map( D => SIG_in(11), CK => clk, Q => n38, 
                           QN => n_2174);
   MY_CLK_r_REG48_S3 : DFF_X1 port map( D => SIG_in(12), CK => clk, Q => n39, 
                           QN => n_2175);
   MY_CLK_r_REG22_S3 : DFF_X1 port map( D => SIG_in(26), CK => clk, Q => n53, 
                           QN => n_2176);
   MY_CLK_r_REG58_S3 : DFF_X2 port map( D => SIG_in(2), CK => clk, Q => n55, QN
                           => n_2177);

end SYN_FPround;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPnormalize_SIG_width28_0 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
         std_logic);

end FPnormalize_SIG_width28_0;

architecture SYN_FPnormalize of FPnormalize_SIG_width28_0 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n7, n9, n11, n12, n14, n15, n17, n32, n33, n34, n35, n36, n37, 
      n38, n39, n40, n41, n42, n43, n44, n45, n46, n48, n49, n50, n51, n52, n53
      , n55, n56, n57, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, 
      n_2190, n_2191, n_2192 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n43, B => n14, ZN => EXP_out(6));
   U9 : NAND3_X1 port map( A1 => n34, A2 => n55, A3 => n33, ZN => n5);
   U11 : XOR2_X1 port map( A => n35, B => n49, Z => EXP_out(2));
   U13 : NOR2_X1 port map( A1 => n48, A2 => n32, ZN => n7);
   U14 : XOR2_X1 port map( A => n37, B => n7, Z => EXP_out(3));
   U15 : NAND3_X1 port map( A1 => n37, A2 => n35, A3 => n49, ZN => n9);
   U16 : INV_X1 port map( A => n9, ZN => n12);
   U17 : XOR2_X1 port map( A => n39, B => n12, Z => EXP_out(4));
   U19 : NOR2_X1 port map( A1 => n50, A2 => n9, ZN => n11);
   U20 : XOR2_X1 port map( A => n41, B => n11, Z => EXP_out(5));
   U21 : NAND3_X1 port map( A1 => n41, A2 => n39, A3 => n12, ZN => n14);
   U23 : NOR2_X1 port map( A1 => n14, A2 => n51, ZN => n15);
   U24 : XOR2_X1 port map( A => n45, B => n15, Z => EXP_out(7));
   U28 : MUX2_X1 port map( A => SIG_in(2), B => SIG_in(3), S => n55, Z => 
                           SIG_out(2));
   U29 : MUX2_X1 port map( A => SIG_in(3), B => SIG_in(4), S => n56, Z => 
                           SIG_out(3));
   U30 : MUX2_X1 port map( A => SIG_in(4), B => SIG_in(5), S => n56, Z => 
                           SIG_out(4));
   U31 : MUX2_X1 port map( A => SIG_in(5), B => SIG_in(6), S => n55, Z => 
                           SIG_out(5));
   U32 : MUX2_X1 port map( A => SIG_in(6), B => SIG_in(7), S => n55, Z => 
                           SIG_out(6));
   U33 : MUX2_X1 port map( A => SIG_in(7), B => SIG_in(8), S => n55, Z => 
                           SIG_out(7));
   U34 : MUX2_X1 port map( A => SIG_in(8), B => SIG_in(9), S => n56, Z => 
                           SIG_out(8));
   U35 : MUX2_X1 port map( A => SIG_in(9), B => SIG_in(10), S => n56, Z => 
                           SIG_out(9));
   U36 : MUX2_X1 port map( A => SIG_in(10), B => SIG_in(11), S => n55, Z => 
                           SIG_out(10));
   U37 : MUX2_X1 port map( A => SIG_in(11), B => SIG_in(12), S => n56, Z => 
                           SIG_out(11));
   U38 : MUX2_X1 port map( A => SIG_in(12), B => SIG_in(13), S => n56, Z => 
                           SIG_out(12));
   U39 : MUX2_X1 port map( A => SIG_in(13), B => SIG_in(14), S => n55, Z => 
                           SIG_out(13));
   U40 : MUX2_X1 port map( A => SIG_in(14), B => SIG_in(15), S => n56, Z => 
                           SIG_out(14));
   U41 : MUX2_X1 port map( A => SIG_in(15), B => SIG_in(16), S => n56, Z => 
                           SIG_out(15));
   U42 : MUX2_X1 port map( A => SIG_in(16), B => SIG_in(17), S => n55, Z => 
                           SIG_out(16));
   U43 : MUX2_X1 port map( A => SIG_in(17), B => SIG_in(18), S => SIG_in(27), Z
                           => SIG_out(17));
   U44 : MUX2_X1 port map( A => SIG_in(18), B => SIG_in(19), S => n56, Z => 
                           SIG_out(18));
   U45 : MUX2_X1 port map( A => SIG_in(19), B => SIG_in(20), S => n55, Z => 
                           SIG_out(19));
   U46 : MUX2_X1 port map( A => SIG_in(20), B => SIG_in(21), S => n55, Z => 
                           SIG_out(20));
   U47 : MUX2_X1 port map( A => SIG_in(21), B => SIG_in(22), S => SIG_in(27), Z
                           => SIG_out(21));
   U48 : MUX2_X1 port map( A => SIG_in(22), B => SIG_in(23), S => n56, Z => 
                           SIG_out(22));
   U49 : MUX2_X1 port map( A => SIG_in(23), B => SIG_in(24), S => n56, Z => 
                           SIG_out(23));
   U50 : MUX2_X1 port map( A => SIG_in(24), B => SIG_in(25), S => n56, Z => 
                           SIG_out(24));
   U51 : MUX2_X1 port map( A => SIG_in(25), B => SIG_in(26), S => n55, Z => 
                           SIG_out(25));
   U52 : INV_X1 port map( A => SIG_in(26), ZN => n17);
   U53 : NAND2_X1 port map( A1 => n17, A2 => n52, ZN => SIG_out(26));
   MY_CLK_r_REG243_S2 : DFF_X1 port map( D => EXP_in(7), CK => clk, Q => n46, 
                           QN => n_2183);
   MY_CLK_r_REG244_S3 : DFF_X1 port map( D => n46, CK => clk, Q => n45, QN => 
                           n_2184);
   MY_CLK_r_REG247_S2 : DFF_X1 port map( D => EXP_in(6), CK => clk, Q => n44, 
                           QN => n_2185);
   MY_CLK_r_REG250_S2 : DFF_X1 port map( D => EXP_in(5), CK => clk, Q => n42, 
                           QN => n_2186);
   MY_CLK_r_REG251_S3 : DFF_X1 port map( D => n42, CK => clk, Q => n41, QN => 
                           n_2187);
   MY_CLK_r_REG253_S2 : DFF_X1 port map( D => EXP_in(4), CK => clk, Q => n40, 
                           QN => n_2188);
   MY_CLK_r_REG256_S2 : DFF_X1 port map( D => EXP_in(3), CK => clk, Q => n38, 
                           QN => n_2189);
   MY_CLK_r_REG257_S3 : DFF_X1 port map( D => n38, CK => clk, Q => n37, QN => 
                           n_2190);
   U4 : INV_X1 port map( A => SIG_in(27), ZN => n52);
   U5 : XNOR2_X1 port map( A => n53, B => n55, ZN => EXP_out(0));
   U6 : CLKBUF_X3 port map( A => SIG_in(27), Z => n55);
   U7 : CLKBUF_X3 port map( A => SIG_in(27), Z => n56);
   U8 : NAND2_X1 port map( A1 => SIG_in(27), A2 => n33, ZN => n57);
   U10 : XNOR2_X1 port map( A => n57, B => n34, ZN => EXP_out(1));
   MY_CLK_r_REG264_S2 : DFF_X1 port map( D => EXP_in(0), CK => clk, Q => n33, 
                           QN => n53);
   MY_CLK_r_REG260_S3 : DFF_X1 port map( D => n36, CK => clk, Q => n35, QN => 
                           n48);
   MY_CLK_r_REG254_S3 : DFF_X1 port map( D => n40, CK => clk, Q => n39, QN => 
                           n50);
   MY_CLK_r_REG248_S3 : DFF_X1 port map( D => n44, CK => clk, Q => n43, QN => 
                           n51);
   MY_CLK_r_REG59_S3 : DFF_X1 port map( D => n5, CK => clk, Q => n32, QN => n49
                           );
   MY_CLK_r_REG262_S2 : DFF_X1 port map( D => EXP_in(1), CK => clk, Q => n34, 
                           QN => n_2191);
   MY_CLK_r_REG259_S2 : DFF_X1 port map( D => EXP_in(2), CK => clk, Q => n36, 
                           QN => n_2192);

end SYN_FPnormalize;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage2_DW01_add_0 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic;  clk : in 
         std_logic);

end FPmul_stage2_DW01_add_0;

architecture SYN_rpl of FPmul_stage2_DW01_add_0 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n2, n_2195, n_2196 : std_logic;

begin
   
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => n2, CO => n_2195, S => 
                           SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1 : OR2_X1 port map( A1 => B(0), A2 => A(0), ZN => carry_1_port);
   U2 : XNOR2_X1 port map( A => B(0), B => A(0), ZN => SUM(0));
   MY_CLK_r_REG245_S1 : DFF_X1 port map( D => carry_7_port, CK => clk, Q => n2,
                           QN => n_2196);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MBE is

   port( A, B : in std_logic_vector (31 downto 0);  C : out std_logic_vector 
         (63 downto 0);  clk : in std_logic);

end MBE;

architecture SYN_beh of MBE is

   component P4_ADDER_NBIT64_NBIT_PER_BLOCK2_NBLOCKS32
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (63 downto 0);  Cout : out std_logic;  clk : 
            in std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_153
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic
            );
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_1
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_2
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_205
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);
   end component;
   
   component FA_206
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co_BAR : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_4
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_5
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_256
      port( A, B, Ci : in std_logic;  Co, S_BAR : out std_logic);
   end component;
   
   component FA_257
      port( A, B, Ci : in std_logic;  Co, S : out std_logic);
   end component;
   
   component FA_258
      port( A, Ci : in std_logic;  Co : out std_logic;  B_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_259
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic
            );
   end component;
   
   component FA_260
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic
            );
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_264
      port( A, B, Ci : in std_logic;  Co, S : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  Co, S : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_268
      port( A, B, Ci : in std_logic;  Co, S : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_7
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_8
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_10
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_11
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_349
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_350
      port( A : in std_logic;  S, Co : out std_logic;  clk, Ci_BAR, B_BAR : in 
            std_logic);
   end component;
   
   component FA_352
      port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_353
      port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_354
      port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_363
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_364
      port( B, Ci : in std_logic;  S, Co : out std_logic;  clk, A_BAR : in 
            std_logic);
   end component;
   
   component FA_365
      port( A, Ci : in std_logic;  S, Co : out std_logic;  clk, B_BAR : in 
            std_logic);
   end component;
   
   component FA_366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_378
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_13
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_14
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_388
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_389
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_390
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_16
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_17
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_19
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_20
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_21
      port( B : in std_logic;  C, S_BAR : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_465
      port( A, B, Ci : in std_logic;  Co : out std_logic;  clk : in std_logic; 
            S_BAR : out std_logic);
   end component;
   
   component FA_466
      port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_476
      port( Ci : in std_logic;  Co : out std_logic;  B_BAR, A_BAR : in 
            std_logic;  S_BAR : out std_logic);
   end component;
   
   component FA_477
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_478
      port( A, B, Ci : in std_logic;  S : out std_logic;  clk : in std_logic;  
            Co_BAR : out std_logic);
   end component;
   
   component FA_479
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_480
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_482
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_22
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_23
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_24
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_485
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_486
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_487
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_488
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_489
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_490
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_491
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_492
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_493
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_25
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_26
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_512
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_513
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_514
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_515
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_516
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_517
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_518
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_519
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_520
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_521
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_522
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_523
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_524
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_525
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_526
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_527
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_528
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_529
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_530
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_531
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_532
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_533
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_534
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_535
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_536
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_28
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_29
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_539
      port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_540
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_541
      port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_542
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_543
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic
            );
   end component;
   
   component FA_544
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_545
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_546
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_547
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_548
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_549
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_550
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_551
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_552
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_553
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_554
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_555
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_556
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_557
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_558
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_559
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_560
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_561
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_562
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_563
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_564
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_565
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_566
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_567
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_568
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_31
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_32
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_33
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_569
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_570
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_571
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_572
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_34
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_35
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_36
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_573
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_574
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_575
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_576
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_577
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_578
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_579
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_580
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_37
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_38
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_39
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_581
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_582
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_583
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_584
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_585
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_586
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_587
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_588
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_589
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_590
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_591
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_592
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_40
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_41
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_42
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_593
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_594
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_595
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_596
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_597
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_598
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_599
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic
            );
   end component;
   
   component FA_600
      port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_601
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_602
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_603
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_604
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_605
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_606
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_607
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_43
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_0
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component ENC_1
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
            p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
            p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
            p_17_port, p_16_port, p_15_port, p_14_BAR, p_13_port, p_12_port, 
            p_11_port, p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, 
            p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, p_0_port : out 
            std_logic);
   end component;
   
   component ENC_2
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
            p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
            p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
            p_17_port, p_16_BAR, p_15_port, p_14_port, p_13_port, p_12_port, 
            p_11_port, p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, 
            p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, p_0_port : out 
            std_logic);
   end component;
   
   component ENC_3
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
            p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
            p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
            p_17_port, p_15_port, p_14_port, p_13_port, p_12_port, p_11_port, 
            p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, p_5_port, 
            p_4_BAR, p_3_port, p_2_port, p_1_port, p_0_port, p_16_BAR : out 
            std_logic);
   end component;
   
   component ENC_4
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
            p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
            p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
            p_17_port, p_15_port, p_14_port, p_13_port, p_12_port, p_11_port, 
            p_10_port, p_9_port, p_8_port, p_7_port, p_6_BAR, p_5_port, 
            p_4_port, p_3_port, p_2_port, p_1_port, p_0_port, p_16_BAR : out 
            std_logic);
   end component;
   
   component ENC_5
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_6
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_7
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_8
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_9
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_10
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_11
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_12
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_13
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_14
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_15
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_16
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_0
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, n207, n208, n209, n210, n211, n212, 
      n213, n214, q_0_0_32_port, q_0_0_31_port, q_0_0_30_port, q_0_0_29_port, 
      q_0_0_28_port, q_0_0_27_port, q_0_0_26_port, q_0_0_25_port, q_0_0_24_port
      , q_0_0_23_port, q_0_0_22_port, q_0_0_21_port, q_0_0_20_port, 
      q_0_0_19_port, q_0_0_18_port, q_0_0_17_port, q_0_0_16_port, q_0_0_15_port
      , q_0_0_14_port, q_0_0_13_port, q_0_0_12_port, q_0_0_11_port, 
      q_0_0_10_port, q_0_0_9_port, q_0_0_8_port, q_0_0_7_port, q_0_0_6_port, 
      q_0_0_5_port, q_0_0_4_port, q_0_0_3_port, q_0_0_2_port, q_0_0_1_port, 
      q_0_0_0_port, q_0_8_47_port, q_0_8_46_port, q_0_8_45_port, q_0_8_44_port,
      q_0_8_43_port, q_0_8_42_port, q_0_8_41_port, q_0_8_40_port, q_0_8_38_port
      , q_0_8_37_port, q_0_8_36_port, q_0_8_35_port, q_0_8_34_port, 
      q_0_8_33_port, q_0_8_32_port, q_0_8_31_port, q_0_8_30_port, q_0_8_29_port
      , q_0_8_28_port, q_0_8_27_port, q_0_8_26_port, q_0_8_25_port, 
      q_0_8_24_port, q_0_8_23_port, q_0_8_22_port, q_0_8_21_port, q_0_8_20_port
      , q_0_8_19_port, q_0_8_18_port, q_0_8_17_port, q_0_8_16_port, 
      q_0_7_47_port, q_0_7_46_port, q_0_7_45_port, q_0_7_44_port, q_0_7_43_port
      , q_0_7_42_port, q_0_7_41_port, q_0_7_40_port, q_0_7_39_port, 
      q_0_7_38_port, q_0_7_37_port, q_0_7_36_port, q_0_7_35_port, q_0_7_34_port
      , q_0_7_33_port, q_0_7_32_port, q_0_7_31_port, q_0_7_30_port, 
      q_0_7_29_port, q_0_7_28_port, q_0_7_27_port, q_0_7_26_port, q_0_7_25_port
      , q_0_7_24_port, q_0_7_23_port, q_0_7_22_port, q_0_7_21_port, 
      q_0_7_20_port, q_0_7_19_port, q_0_7_18_port, q_0_7_17_port, q_0_7_16_port
      , q_0_7_15_port, q_0_7_14_port, q_0_6_47_port, q_0_6_46_port, 
      q_0_6_45_port, q_0_6_44_port, q_0_6_43_port, q_0_6_42_port, q_0_6_41_port
      , q_0_6_40_port, q_0_6_39_port, q_0_6_38_port, q_0_6_37_port, 
      q_0_6_36_port, q_0_6_35_port, q_0_6_34_port, q_0_6_33_port, q_0_6_32_port
      , q_0_6_31_port, q_0_6_30_port, q_0_6_29_port, q_0_6_28_port, 
      q_0_6_27_port, q_0_6_26_port, q_0_6_25_port, q_0_6_24_port, q_0_6_23_port
      , q_0_6_22_port, q_0_6_21_port, q_0_6_20_port, q_0_6_19_port, 
      q_0_6_18_port, q_0_6_17_port, q_0_6_16_port, q_0_6_15_port, q_0_6_14_port
      , q_0_6_13_port, q_0_6_12_port, q_0_5_47_port, q_0_5_46_port, 
      q_0_5_45_port, q_0_5_44_port, q_0_5_43_port, q_0_5_42_port, q_0_5_41_port
      , q_0_5_40_port, q_0_5_39_port, q_0_5_38_port, q_0_5_37_port, 
      q_0_5_36_port, q_0_5_35_port, q_0_5_34_port, q_0_5_33_port, q_0_5_32_port
      , q_0_5_31_port, q_0_5_30_port, q_0_5_29_port, q_0_5_28_port, 
      q_0_5_27_port, q_0_5_26_port, q_0_5_25_port, q_0_5_24_port, q_0_5_23_port
      , q_0_5_22_port, q_0_5_21_port, q_0_5_20_port, q_0_5_19_port, 
      q_0_5_18_port, q_0_5_17_port, q_0_5_16_port, q_0_5_15_port, q_0_5_14_port
      , q_0_5_13_port, q_0_5_12_port, q_0_5_11_port, q_0_5_10_port, 
      q_0_4_47_port, q_0_4_46_port, q_0_4_45_port, q_0_4_44_port, q_0_4_43_port
      , q_0_4_42_port, q_0_4_41_port, q_0_4_40_port, q_0_4_39_port, 
      q_0_4_38_port, q_0_4_37_port, q_0_4_36_port, q_0_4_35_port, q_0_4_34_port
      , q_0_4_33_port, q_0_4_32_port, q_0_4_31_port, q_0_4_30_port, 
      q_0_4_29_port, q_0_4_28_port, q_0_4_27_port, q_0_4_26_port, q_0_4_25_port
      , q_0_4_24_port, q_0_4_23_port, q_0_4_22_port, q_0_4_21_port, 
      q_0_4_20_port, q_0_4_19_port, q_0_4_18_port, q_0_4_17_port, q_0_4_16_port
      , q_0_4_15_port, q_0_4_14_port, q_0_4_13_port, q_0_4_12_port, 
      q_0_4_11_port, q_0_4_10_port, q_0_4_9_port, q_0_4_8_port, q_0_3_47_port, 
      q_0_3_46_port, q_0_3_45_port, q_0_3_44_port, q_0_3_43_port, q_0_3_42_port
      , q_0_3_41_port, q_0_3_40_port, q_0_3_39_port, q_0_3_38_port, 
      q_0_3_37_port, q_0_3_36_port, q_0_3_35_port, q_0_3_34_port, q_0_3_33_port
      , q_0_3_32_port, q_0_3_31_port, q_0_3_30_port, q_0_3_29_port, 
      q_0_3_28_port, q_0_3_27_port, q_0_3_26_port, q_0_3_25_port, q_0_3_24_port
      , q_0_3_23_port, q_0_3_22_port, q_0_3_21_port, q_0_3_20_port, 
      q_0_3_19_port, q_0_3_18_port, q_0_3_17_port, q_0_3_16_port, q_0_3_15_port
      , q_0_3_14_port, q_0_3_13_port, q_0_3_12_port, q_0_3_11_port, 
      q_0_3_10_port, q_0_3_9_port, q_0_3_8_port, q_0_3_7_port, q_0_3_6_port, 
      q_0_2_47_port, q_0_2_46_port, q_0_2_45_port, q_0_2_44_port, q_0_2_43_port
      , q_0_2_42_port, q_0_2_41_port, q_0_2_40_port, q_0_2_39_port, 
      q_0_2_38_port, q_0_2_37_port, q_0_2_36_port, q_0_2_35_port, q_0_2_34_port
      , q_0_2_33_port, q_0_2_32_port, q_0_2_31_port, q_0_2_30_port, 
      q_0_2_29_port, q_0_2_28_port, q_0_2_27_port, q_0_2_26_port, q_0_2_25_port
      , q_0_2_24_port, q_0_2_23_port, q_0_2_22_port, q_0_2_21_port, 
      q_0_2_20_port, q_0_2_19_port, q_0_2_18_port, q_0_2_17_port, q_0_2_16_port
      , q_0_2_15_port, q_0_2_14_port, q_0_2_13_port, q_0_2_12_port, 
      q_0_2_11_port, q_0_2_10_port, q_0_2_9_port, q_0_2_8_port, q_0_2_7_port, 
      q_0_2_6_port, q_0_2_5_port, q_0_2_4_port, q_0_1_47_port, q_0_1_46_port, 
      q_0_1_45_port, q_0_1_44_port, q_0_1_43_port, q_0_1_42_port, q_0_1_41_port
      , q_0_1_40_port, q_0_1_39_port, q_0_1_38_port, q_0_1_37_port, 
      q_0_1_36_port, q_0_1_34_port, q_0_1_33_port, q_0_1_32_port, q_0_1_31_port
      , q_0_1_30_port, q_0_1_29_port, q_0_1_28_port, q_0_1_27_port, 
      q_0_1_26_port, q_0_1_25_port, q_0_1_24_port, q_0_1_23_port, q_0_1_22_port
      , q_0_1_21_port, q_0_1_20_port, q_0_1_19_port, q_0_1_18_port, 
      q_0_1_17_port, q_0_1_16_port, q_0_1_15_port, q_0_1_14_port, q_0_1_13_port
      , q_0_1_12_port, q_0_1_11_port, q_0_1_10_port, q_0_1_9_port, q_0_1_8_port
      , q_0_1_7_port, q_0_1_6_port, q_0_1_5_port, q_0_1_4_port, q_0_1_3_port, 
      q_0_1_2_port, q_0_14_32_port, q_0_14_31_port, q_0_14_30_port, 
      q_0_14_29_port, q_0_14_28_port, q_0_13_32_port, q_0_13_31_port, 
      q_0_13_30_port, q_0_13_29_port, q_0_13_28_port, q_0_13_27_port, 
      q_0_13_26_port, q_0_12_35_port, q_0_12_34_port, q_0_12_33_port, 
      q_0_12_32_port, q_0_12_31_port, q_0_12_30_port, q_0_12_29_port, 
      q_0_12_28_port, q_0_12_27_port, q_0_12_26_port, q_0_12_25_port, 
      q_0_12_24_port, q_0_11_36_port, q_0_11_35_port, q_0_11_34_port, 
      q_0_11_33_port, q_0_11_32_port, q_0_11_31_port, q_0_11_30_port, 
      q_0_11_29_port, q_0_11_28_port, q_0_11_27_port, q_0_11_26_port, 
      q_0_11_25_port, q_0_11_24_port, q_0_11_23_port, q_0_11_22_port, 
      q_0_10_46_port, q_0_10_38_port, q_0_10_37_port, q_0_10_36_port, 
      q_0_10_35_port, q_0_10_34_port, q_0_10_33_port, q_0_10_32_port, 
      q_0_10_31_port, q_0_10_30_port, q_0_10_29_port, q_0_10_28_port, 
      q_0_10_27_port, q_0_10_26_port, q_0_10_25_port, q_0_10_24_port, 
      q_0_10_23_port, q_0_10_22_port, q_0_10_21_port, q_0_10_20_port, 
      q_0_9_47_port, q_0_9_46_port, q_0_9_44_port, q_0_9_42_port, q_0_9_40_port
      , q_0_9_39_port, q_0_9_38_port, q_0_9_37_port, q_0_9_36_port, 
      q_0_9_35_port, q_0_9_34_port, q_0_9_33_port, q_0_9_32_port, q_0_9_31_port
      , q_0_9_30_port, q_0_9_29_port, q_0_9_28_port, q_0_9_27_port, 
      q_0_9_26_port, q_0_9_25_port, q_0_9_24_port, q_0_9_23_port, q_0_9_22_port
      , q_0_9_21_port, q_0_9_20_port, q_0_9_19_port, q_0_9_18_port, 
      q_1_1_42_port, q_1_1_41_port, q_1_1_40_port, q_1_1_39_port, q_1_1_38_port
      , q_1_1_37_port, q_1_1_36_port, q_1_1_35_port, q_1_1_34_port, 
      q_1_1_33_port, q_1_1_32_port, q_1_1_31_port, q_1_1_30_port, q_1_1_29_port
      , q_1_1_28_port, q_1_1_27_port, q_1_1_26_port, q_1_1_25_port, 
      q_1_0_43_port, q_1_0_42_port, q_1_0_41_port, q_1_0_40_port, q_1_0_39_port
      , q_1_0_38_port, q_1_0_37_port, q_1_0_36_port, q_1_0_35_port, 
      q_1_0_34_port, q_1_0_33_port, q_1_0_32_port, q_1_0_31_port, q_1_0_30_port
      , q_1_0_29_port, q_1_0_28_port, q_1_0_27_port, q_1_0_26_port, 
      q_1_0_25_port, q_1_0_24_port, q_1_7_35_port, q_1_7_34_port, q_1_7_33_port
      , q_1_7_32_port, q_1_7_31_port, q_1_6_37_port, q_1_6_36_port, 
      q_1_6_35_port, q_1_6_34_port, q_1_6_33_port, q_1_6_32_port, q_1_6_31_port
      , q_1_5_38_port, q_1_5_37_port, q_1_5_36_port, q_1_5_34_port, 
      q_1_5_33_port, q_1_5_32_port, q_1_5_31_port, q_1_5_30_port, q_1_5_29_port
      , q_1_4_39_port, q_1_4_38_port, q_1_4_37_port, q_1_4_36_port, 
      q_1_4_35_port, q_1_4_34_port, q_1_4_33_port, q_1_4_32_port, q_1_4_31_port
      , q_1_4_30_port, q_1_4_29_port, q_1_4_28_port, q_1_3_40_port, 
      q_1_3_39_port, q_1_3_38_port, q_1_3_37_port, q_1_3_36_port, q_1_3_35_port
      , q_1_3_34_port, q_1_3_33_port, q_1_3_32_port, q_1_3_31_port, 
      q_1_3_29_port, q_1_3_28_port, q_1_3_27_port, q_1_2_41_port, q_1_2_40_port
      , q_1_2_39_port, q_1_2_38_port, q_1_2_37_port, q_1_2_35_port, 
      q_1_2_34_port, q_1_2_33_port, q_1_2_32_port, q_1_2_30_port, q_1_2_29_port
      , q_1_2_28_port, q_1_2_27_port, q_1_2_26_port, q_2_2_47_port, 
      q_2_2_46_port, q_2_2_45_port, q_2_2_44_port, q_2_2_43_port, q_2_2_42_port
      , q_2_2_41_port, q_2_2_40_port, q_2_2_39_port, q_2_2_38_port, 
      q_2_2_37_port, q_2_2_36_port, q_2_2_35_port, q_2_2_34_port, q_2_2_33_port
      , q_2_2_32_port, q_2_2_31_port, q_2_2_30_port, q_2_2_29_port, 
      q_2_2_28_port, q_2_2_27_port, q_2_2_26_port, q_2_2_25_port, q_2_2_23_port
      , q_2_2_22_port, q_2_2_21_port, q_2_2_20_port, q_2_2_19_port, 
      q_2_2_18_port, q_2_1_47_port, q_2_1_46_port, q_2_1_45_port, q_2_1_44_port
      , q_2_1_43_port, q_2_1_42_port, q_2_1_41_port, q_2_1_40_port, 
      q_2_1_39_port, q_2_1_38_port, q_2_1_37_port, q_2_1_36_port, q_2_1_35_port
      , q_2_1_34_port, q_2_1_33_port, q_2_1_32_port, q_2_1_31_port, 
      q_2_1_30_port, q_2_1_29_port, q_2_1_28_port, q_2_1_27_port, q_2_1_26_port
      , q_2_1_25_port, q_2_1_24_port, q_2_1_23_port, q_2_1_22_port, 
      q_2_1_21_port, q_2_1_20_port, q_2_1_19_port, q_2_1_18_port, q_2_1_17_port
      , q_2_0_47_port, q_2_0_46_port, q_2_0_45_port, q_2_0_44_port, 
      q_2_0_43_port, q_2_0_42_port, q_2_0_41_port, q_2_0_40_port, q_2_0_39_port
      , q_2_0_38_port, q_2_0_37_port, q_2_0_36_port, q_2_0_35_port, 
      q_2_0_34_port, q_2_0_33_port, q_2_0_32_port, q_2_0_31_port, q_2_0_30_port
      , q_2_0_29_port, q_2_0_28_port, q_2_0_27_port, q_2_0_26_port, 
      q_2_0_25_port, q_2_0_24_port, q_2_0_23_port, q_2_0_22_port, q_2_0_21_port
      , q_2_0_20_port, q_2_0_19_port, q_2_0_18_port, q_2_0_17_port, 
      q_2_0_16_port, q_2_7_33_port, q_2_7_32_port, q_2_7_31_port, q_2_7_30_port
      , q_2_7_29_port, q_2_7_28_port, q_2_7_27_port, q_2_7_26_port, 
      q_2_7_25_port, q_2_7_24_port, q_2_7_23_port, q_2_6_44_port, q_2_6_43_port
      , q_2_6_42_port, q_2_6_32_port, q_2_6_31_port, q_2_6_30_port, 
      q_2_6_28_port, q_2_6_27_port, q_2_6_26_port, q_2_6_25_port, q_2_6_24_port
      , q_2_6_23_port, q_2_6_22_port, q_2_5_46_port, q_2_5_45_port, 
      q_2_5_44_port, q_2_5_43_port, q_2_5_42_port, q_2_5_41_port, q_2_5_40_port
      , q_2_5_39_port, q_2_5_38_port, q_2_5_37_port, q_2_5_36_port, 
      q_2_5_35_port, q_2_5_34_port, q_2_5_33_port, q_2_5_32_port, q_2_5_31_port
      , q_2_5_30_port, q_2_5_29_port, q_2_5_28_port, q_2_5_27_port, 
      q_2_5_26_port, q_2_5_25_port, q_2_5_24_port, q_2_5_23_port, q_2_5_22_port
      , q_2_5_21_port, q_2_4_47_port, q_2_4_46_port, q_2_4_45_port, 
      q_2_4_44_port, q_2_4_43_port, q_2_4_42_port, q_2_4_41_port, q_2_4_40_port
      , q_2_4_39_port, q_2_4_38_port, q_2_4_37_port, q_2_4_36_port, 
      q_2_4_35_port, q_2_4_34_port, q_2_4_33_port, q_2_4_32_port, q_2_4_31_port
      , q_2_4_30_port, q_2_4_29_port, q_2_4_28_port, q_2_4_27_port, 
      q_2_4_26_port, q_2_4_25_port, q_2_4_24_port, q_2_4_23_port, q_2_4_22_port
      , q_2_3_47_port, q_2_3_46_port, q_2_3_45_port, q_2_3_44_port, 
      q_2_3_43_port, q_2_3_42_port, q_2_3_41_port, q_2_3_40_port, q_2_3_39_port
      , q_2_3_38_port, q_2_3_37_port, q_2_3_36_port, q_2_3_35_port, 
      q_2_3_34_port, q_2_3_33_port, q_2_3_32_port, q_2_3_31_port, q_2_3_30_port
      , q_2_3_29_port, q_2_3_28_port, q_2_3_27_port, q_2_3_26_port, 
      q_2_3_25_port, q_2_3_24_port, q_2_3_23_port, q_2_3_22_port, q_2_3_21_port
      , q_2_3_20_port, q_2_3_19_port, q_3_3_47_port, q_3_3_46_port, 
      q_3_3_45_port, q_3_3_44_port, q_3_3_43_port, q_3_3_42_port, q_3_3_41_port
      , q_3_3_40_port, q_3_3_39_port, q_3_3_38_port, q_3_3_37_port, 
      q_3_3_36_port, q_3_3_35_port, q_3_3_34_port, q_3_3_33_port, q_3_3_32_port
      , q_3_3_31_port, q_3_3_30_port, q_3_3_29_port, q_3_3_28_port, 
      q_3_3_27_port, q_3_3_26_port, q_3_3_25_port, q_3_3_24_port, q_3_3_23_port
      , q_3_3_22_port, q_3_3_21_port, q_3_3_20_port, q_3_3_19_port, 
      q_3_3_18_port, q_3_3_17_port, q_3_3_16_port, q_3_3_15_port, q_3_3_14_port
      , q_3_3_13_port, q_3_2_47_port, q_3_2_46_port, q_3_2_45_port, 
      q_3_2_44_port, q_3_2_43_port, q_3_2_42_port, q_3_2_41_port, q_3_2_40_port
      , q_3_2_39_port, q_3_2_38_port, q_3_2_37_port, q_3_2_36_port, 
      q_3_2_35_port, q_3_2_34_port, q_3_2_33_port, q_3_2_32_port, q_3_2_31_port
      , q_3_2_30_port, q_3_2_29_port, q_3_2_28_port, q_3_2_27_port, 
      q_3_2_26_port, q_3_2_25_port, q_3_2_24_port, q_3_2_23_port, q_3_2_22_port
      , q_3_2_21_port, q_3_2_20_port, q_3_2_19_port, q_3_2_18_port, 
      q_3_2_17_port, q_3_2_16_port, q_3_2_15_port, q_3_2_14_port, q_3_2_13_port
      , q_3_2_12_port, q_3_1_47_port, q_3_1_46_port, q_3_1_45_port, 
      q_3_1_44_port, q_3_1_43_port, q_3_1_42_port, q_3_1_41_port, q_3_1_40_port
      , q_3_1_39_port, q_3_1_38_port, q_3_1_37_port, q_3_1_36_port, 
      q_3_1_35_port, q_3_1_34_port, q_3_1_33_port, q_3_1_32_port, q_3_1_31_port
      , q_3_1_30_port, q_3_1_29_port, q_3_1_28_port, q_3_1_27_port, 
      q_3_1_26_port, q_3_1_25_port, q_3_1_24_port, q_3_1_23_port, q_3_1_22_port
      , q_3_1_21_port, q_3_1_20_port, q_3_1_19_port, q_3_1_18_port, 
      q_3_1_17_port, q_3_1_16_port, q_3_1_15_port, q_3_1_14_port, q_3_1_13_port
      , q_3_1_12_port, q_3_1_11_port, q_3_0_47_port, q_3_0_46_port, 
      q_3_0_45_port, q_3_0_44_port, q_3_0_43_port, q_3_0_42_port, q_3_0_41_port
      , q_3_0_40_port, q_3_0_39_port, q_3_0_38_port, q_3_0_37_port, 
      q_3_0_36_port, q_3_0_35_port, q_3_0_34_port, q_3_0_33_port, q_3_0_32_port
      , q_3_0_31_port, q_3_0_30_port, q_3_0_29_port, q_3_0_28_port, 
      q_3_0_25_port, q_3_0_24_port, q_3_0_23_port, q_3_0_22_port, q_3_0_21_port
      , q_3_0_20_port, q_3_0_19_port, q_3_0_18_port, q_3_0_17_port, 
      q_3_0_16_port, q_3_0_15_port, q_3_0_14_port, q_3_0_13_port, q_3_0_11_port
      , q_3_5_47_port, q_3_5_33_port, q_3_5_32_port, q_3_5_31_port, 
      q_3_5_30_port, q_3_5_29_port, q_3_5_28_port, q_3_5_27_port, q_3_5_26_port
      , q_3_5_25_port, q_3_5_24_port, q_3_5_23_port, q_3_5_22_port, 
      q_3_5_21_port, q_3_5_20_port, q_3_5_19_port, q_3_5_18_port, q_3_5_17_port
      , q_3_5_16_port, q_3_5_15_port, q_3_4_47_port, q_3_4_46_port, 
      q_3_4_44_port, q_3_4_43_port, q_3_4_42_port, q_3_4_33_port, q_3_4_32_port
      , q_3_4_31_port, q_3_4_30_port, q_3_4_29_port, q_3_4_28_port, 
      q_3_4_27_port, q_3_4_26_port, q_3_4_25_port, q_3_4_24_port, q_3_4_23_port
      , q_3_4_22_port, q_3_4_21_port, q_3_4_20_port, q_3_4_19_port, 
      q_3_4_18_port, q_3_4_17_port, q_3_4_16_port, q_3_4_15_port, q_4_2_47_port
      , q_4_2_46_port, q_4_2_45_port, q_4_2_44_port, q_4_2_43_port, 
      q_4_2_42_port, q_4_2_41_port, q_4_2_40_port, q_4_2_39_port, q_4_2_38_port
      , q_4_2_37_port, q_4_2_36_port, q_4_2_35_port, q_4_2_34_port, 
      q_4_2_33_port, q_4_2_32_port, q_4_2_31_port, q_4_2_30_port, q_4_2_29_port
      , q_4_2_28_port, q_4_2_27_port, q_4_2_26_port, q_4_2_25_port, 
      q_4_2_24_port, q_4_2_21_port, q_4_2_19_port, q_4_2_18_port, q_4_2_17_port
      , q_4_2_16_port, q_4_2_15_port, q_4_2_14_port, q_4_2_13_port, 
      q_4_2_12_port, q_4_2_11_port, q_4_2_10_port, q_4_2_9_port, q_4_2_8_port, 
      q_4_1_47_port, q_4_1_46_port, q_4_1_45_port, q_4_1_44_port, q_4_1_43_port
      , q_4_1_42_port, q_4_1_41_port, q_4_1_40_port, q_4_1_39_port, 
      q_4_1_38_port, q_4_1_37_port, q_4_1_36_port, q_4_1_35_port, q_4_1_34_port
      , q_4_1_33_port, q_4_1_32_port, q_4_1_31_port, q_4_1_30_port, 
      q_4_1_29_port, q_4_1_28_port, q_4_1_27_port, q_4_1_26_port, q_4_1_25_port
      , q_4_1_24_port, q_4_1_23_port, q_4_1_22_port, q_4_1_21_port, 
      q_4_1_20_port, q_4_1_19_port, q_4_1_18_port, q_4_1_17_port, q_4_1_16_port
      , q_4_1_15_port, q_4_1_14_port, q_4_1_13_port, q_4_1_12_port, 
      q_4_1_11_port, q_4_1_10_port, q_4_1_9_port, q_4_1_8_port, q_4_1_7_port, 
      q_4_0_47_port, q_4_0_46_port, q_4_0_45_port, q_4_0_44_port, q_4_0_43_port
      , q_4_0_42_port, q_4_0_41_port, q_4_0_40_port, q_4_0_39_port, 
      q_4_0_38_port, q_4_0_37_port, q_4_0_36_port, q_4_0_35_port, q_4_0_34_port
      , q_4_0_33_port, q_4_0_32_port, q_4_0_31_port, q_4_0_30_port, 
      q_4_0_29_port, q_4_0_28_port, q_4_0_27_port, q_4_0_26_port, q_4_0_24_port
      , q_4_0_21_port, q_4_0_20_port, q_4_0_19_port, q_4_0_18_port, 
      q_4_0_17_port, q_4_0_16_port, q_4_0_15_port, q_4_0_14_port, q_4_0_13_port
      , q_4_0_12_port, q_4_0_11_port, q_4_0_10_port, q_4_0_9_port, q_4_0_8_port
      , q_4_0_7_port, q_4_0_6_port, q_5_2_47_port, q_5_2_45_port, q_5_2_44_port
      , q_5_2_43_port, q_5_2_34_port, q_5_2_33_port, q_5_2_32_port, 
      q_5_2_31_port, q_5_2_30_port, q_5_2_29_port, q_5_2_28_port, q_5_2_27_port
      , q_5_2_26_port, q_5_2_25_port, q_5_2_24_port, q_5_2_23_port, 
      q_5_2_22_port, q_5_2_21_port, q_5_2_20_port, q_5_2_19_port, q_5_2_18_port
      , q_5_2_17_port, q_5_2_16_port, q_5_2_15_port, q_5_2_14_port, 
      q_5_2_13_port, q_5_2_12_port, q_5_2_11_port, q_5_2_10_port, q_5_2_9_port,
      q_5_1_47_port, q_5_1_46_port, q_5_1_45_port, q_5_1_44_port, q_5_1_43_port
      , q_5_1_42_port, q_5_1_41_port, q_5_1_40_port, q_5_1_39_port, 
      q_5_1_38_port, q_5_1_37_port, q_5_1_36_port, q_5_1_35_port, q_5_1_34_port
      , q_5_1_33_port, q_5_1_32_port, q_5_1_31_port, q_5_1_30_port, 
      q_5_1_29_port, q_5_1_28_port, q_5_1_27_port, q_5_1_26_port, q_5_1_25_port
      , q_5_1_24_port, q_5_1_23_port, q_5_1_22_port, q_5_1_21_port, 
      q_5_1_20_port, q_5_1_19_port, q_5_1_18_port, q_5_1_17_port, q_5_1_16_port
      , q_5_1_15_port, q_5_1_14_port, q_5_1_13_port, q_5_1_12_port, 
      q_5_1_11_port, q_5_1_10_port, q_5_1_9_port, q_5_1_8_port, q_5_1_7_port, 
      q_5_1_6_port, q_5_1_5_port, q_5_0_47_port, q_5_0_46_port, q_5_0_45_port, 
      q_5_0_44_port, q_5_0_43_port, q_5_0_42_port, q_5_0_41_port, q_5_0_40_port
      , q_5_0_39_port, q_5_0_38_port, q_5_0_37_port, q_5_0_36_port, 
      q_5_0_35_port, q_5_0_34_port, q_5_0_33_port, q_5_0_32_port, q_5_0_31_port
      , q_5_0_30_port, q_5_0_29_port, q_5_0_28_port, q_5_0_27_port, 
      q_5_0_26_port, q_5_0_25_port, q_5_0_24_port, q_5_0_23_port, q_5_0_22_port
      , q_5_0_21_port, q_5_0_20_port, q_5_0_19_port, q_5_0_18_port, 
      q_5_0_17_port, q_5_0_15_port, q_5_0_14_port, q_5_0_13_port, q_5_0_12_port
      , q_5_0_11_port, q_5_0_10_port, q_5_0_9_port, q_5_0_8_port, q_5_0_7_port,
      q_5_0_6_port, q_5_0_5_port, q_5_0_4_port, q_6_1_47_port, q_6_1_46_port, 
      q_6_1_45_port, q_6_1_44_port, q_6_1_43_port, q_6_1_42_port, q_6_1_41_port
      , q_6_1_40_port, q_6_1_39_port, q_6_1_38_port, q_6_1_37_port, 
      q_6_1_36_port, q_6_1_34_port, q_6_1_32_port, q_6_1_31_port, q_6_1_30_port
      , q_6_1_28_port, q_6_1_26_port, q_6_1_25_port, q_6_1_24_port, 
      q_6_1_23_port, q_6_1_22_port, q_6_1_21_port, q_6_1_20_port, q_6_1_19_port
      , q_6_1_18_port, q_6_1_17_port, q_6_1_16_port, q_6_1_15_port, 
      q_6_1_14_port, q_6_1_13_port, q_6_1_12_port, q_6_1_11_port, q_6_1_10_port
      , q_6_1_9_port, q_6_1_8_port, q_6_1_7_port, q_6_1_6_port, q_6_1_5_port, 
      q_6_1_4_port, q_6_1_3_port, q_6_0_47_port, q_6_0_46_port, q_6_0_45_port, 
      q_6_0_44_port, q_6_0_43_port, q_6_0_42_port, q_6_0_41_port, q_6_0_40_port
      , q_6_0_38_port, q_6_0_37_port, q_6_0_36_port, q_6_0_35_port, 
      q_6_0_34_port, q_6_0_32_port, q_6_0_31_port, q_6_0_30_port, q_6_0_29_port
      , q_6_0_28_port, q_6_0_27_port, q_6_0_26_port, q_6_0_25_port, 
      q_6_0_24_port, q_6_0_23_port, q_6_0_22_port, q_6_0_21_port, q_6_0_20_port
      , q_6_0_19_port, q_6_0_18_port, q_6_0_17_port, q_6_0_16_port, 
      q_6_0_15_port, q_6_0_14_port, q_6_0_13_port, q_6_0_12_port, q_6_0_11_port
      , q_6_0_10_port, q_6_0_9_port, q_6_0_8_port, q_6_0_7_port, q_6_0_6_port, 
      q_6_0_5_port, q_6_0_4_port, q_6_0_3_port, q_6_0_2_port, n2, n91, n92, n93
      , n95, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n205, 
      net102724, net102725, net102726, net102727, net102728, net102729, 
      net102730, net102731, net102732, net102733, net102734, net102735, 
      net102736, net102737, net102738, net102739, net102740, net102741, 
      net102742, net102743, net102744, net102745, net102746, net102747, 
      net102748, net102749, net102750, net102751, net102752, net102753, 
      net102754, net102755, net102756, net102757, net102758, net102759, 
      net102760, net102761, net102762, net102763, net102764, net102765, 
      net102766, net102767, net102768, net102769, net102770, net102771, 
      net102772, net102773, net102774, net102775, net102776, net102777, 
      net102778, net102779, net102780, net102781, net102782, net102783, 
      net102784, net102785, net102786, net102787, net102788, net102789, 
      net102790, net102791, net102792, net102793, net102794, net102795, 
      net102796, net102797, net102798, net102799, net102800, net102801, 
      net102802, net102803, net102804, net102805, net102806, net102807, 
      net102808, net102809, net102810, net102811, net102812, net102813, 
      net102814, net102815, net102816, net102817, net102818, net102819, 
      net102820, net102821, net102822, net102823, n_2251, n_2252, n_2253, 
      n_2254, n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, 
      n_2263, n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, 
      n_2272, n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, 
      n_2281, n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, 
      n_2290, n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, 
      n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, 
      n_2308, n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, 
      n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, 
      n_2326, n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, 
      n_2335, n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, 
      n_2344, n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, 
      n_2353, n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, 
      n_2362, n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, 
      n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, 
      n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, 
      n_2389, n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, 
      n_2398, n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, 
      n_2407, n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, 
      n_2416, n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, 
      n_2425, n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, 
      n_2434, n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, 
      n_2443, n_2444, n_2445 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   U4 : CLKBUF_X1 port map( A => B(23), Z => n2);
   U93 : INV_X1 port map( A => B(9), ZN => n91);
   U94 : INV_X1 port map( A => B(7), ZN => n92);
   U95 : INV_X1 port map( A => B(5), ZN => n93);
   U97 : INV_X1 port map( A => B(1), ZN => n95);
   n120 <= '0';
   n121 <= '0';
   n122 <= '0';
   n123 <= '0';
   n124 <= '0';
   n125 <= '0';
   n126 <= '0';
   n127 <= '0';
   n128 <= '0';
   n129 <= '0';
   n130 <= '0';
   n131 <= '0';
   n132 <= '0';
   n133 <= '0';
   n134 <= '0';
   n135 <= '0';
   n136 <= '0';
   n137 <= '0';
   n138 <= '0';
   n139 <= '0';
   n140 <= '0';
   n141 <= '0';
   n142 <= '0';
   n143 <= '0';
   n144 <= '0';
   n145 <= '0';
   n146 <= '0';
   n147 <= '0';
   n148 <= '0';
   n149 <= '0';
   n150 <= '0';
   n151 <= '0';
   n152 <= '0';
   n153 <= '0';
   n154 <= '0';
   n155 <= '0';
   n156 <= '0';
   n157 <= '0';
   n158 <= '0';
   n159 <= '0';
   n160 <= '0';
   n161 <= '0';
   n162 <= '0';
   n163 <= '0';
   n164 <= '0';
   n165 <= '0';
   n166 <= '0';
   n167 <= '0';
   n168 <= '0';
   n169 <= '0';
   n170 <= '0';
   n171 <= '0';
   n214 <= '0';
   n213 <= '0';
   n212 <= '0';
   n211 <= '0';
   n210 <= '0';
   n209 <= '0';
   n208 <= '0';
   n207 <= '0';
   n205 <= '0';
   net102724 <= '0';
   net102725 <= '0';
   net102726 <= '0';
   net102727 <= '0';
   net102728 <= '0';
   net102729 <= '0';
   net102730 <= '0';
   net102731 <= '0';
   net102732 <= '0';
   net102733 <= '0';
   net102734 <= '0';
   net102735 <= '0';
   net102736 <= '0';
   net102737 <= '0';
   net102738 <= '0';
   net102739 <= '0';
   net102740 <= '0';
   net102741 <= '0';
   net102742 <= '0';
   net102743 <= '0';
   net102744 <= '0';
   net102745 <= '0';
   net102746 <= '0';
   net102747 <= '0';
   net102748 <= '0';
   net102749 <= '0';
   net102750 <= '0';
   net102751 <= '0';
   net102752 <= '0';
   net102753 <= '0';
   net102754 <= '0';
   net102755 <= '0';
   net102756 <= '0';
   net102757 <= '0';
   net102758 <= '0';
   net102759 <= '0';
   net102760 <= '0';
   net102761 <= '0';
   net102762 <= '0';
   net102763 <= '0';
   net102764 <= '0';
   net102765 <= '0';
   net102766 <= '0';
   net102767 <= '0';
   net102768 <= '0';
   net102769 <= '0';
   net102770 <= '0';
   net102771 <= '0';
   net102772 <= '0';
   net102773 <= '0';
   net102774 <= '0';
   net102775 <= '0';
   net102776 <= '0';
   net102777 <= '0';
   net102778 <= '0';
   net102779 <= '0';
   net102780 <= '0';
   net102781 <= '0';
   net102782 <= '0';
   net102783 <= '0';
   net102784 <= '0';
   net102785 <= '0';
   net102786 <= '0';
   net102787 <= '0';
   net102788 <= '0';
   net102789 <= '0';
   net102790 <= '0';
   net102791 <= '0';
   net102792 <= '0';
   net102793 <= '0';
   net102794 <= '0';
   net102795 <= '0';
   net102796 <= '0';
   net102797 <= '0';
   net102798 <= '0';
   net102799 <= '0';
   net102800 <= '0';
   net102801 <= '0';
   net102802 <= '0';
   net102803 <= '0';
   net102804 <= '0';
   net102805 <= '0';
   net102806 <= '0';
   net102807 <= '0';
   net102808 <= '0';
   net102809 <= '0';
   net102810 <= '0';
   net102811 <= '0';
   net102812 <= '0';
   net102813 <= '0';
   net102814 <= '0';
   net102815 <= '0';
   net102816 <= '0';
   net102817 <= '0';
   net102818 <= '0';
   net102819 <= '0';
   net102820 <= '0';
   net102821 <= '0';
   net102822 <= '0';
   net102823 <= '0';
   encI_1 : ENC_0 port map( b(2) => B(1), b(1) => B(0), b(0) => X_Logic0_port, 
                           A(31) => n205, A(30) => n205, A(29) => n205, A(28) 
                           => n205, A(27) => n205, A(26) => n205, A(25) => n205
                           , A(24) => n205, A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), p(32) => 
                           q_0_0_32_port, p(31) => q_0_0_31_port, p(30) => 
                           q_0_0_30_port, p(29) => q_0_0_29_port, p(28) => 
                           q_0_0_28_port, p(27) => q_0_0_27_port, p(26) => 
                           q_0_0_26_port, p(25) => q_0_0_25_port, p(24) => 
                           q_0_0_24_port, p(23) => q_0_0_23_port, p(22) => 
                           q_0_0_22_port, p(21) => q_0_0_21_port, p(20) => 
                           q_0_0_20_port, p(19) => q_0_0_19_port, p(18) => 
                           q_0_0_18_port, p(17) => q_0_0_17_port, p(16) => 
                           q_0_0_16_port, p(15) => q_0_0_15_port, p(14) => 
                           q_0_0_14_port, p(13) => q_0_0_13_port, p(12) => 
                           q_0_0_12_port, p(11) => q_0_0_11_port, p(10) => 
                           q_0_0_10_port, p(9) => q_0_0_9_port, p(8) => 
                           q_0_0_8_port, p(7) => q_0_0_7_port, p(6) => 
                           q_0_0_6_port, p(5) => q_0_0_5_port, p(4) => 
                           q_0_0_4_port, p(3) => q_0_0_3_port, p(2) => 
                           q_0_0_2_port, p(1) => q_0_0_1_port, p(0) => 
                           q_0_0_0_port);
   encI_2 : ENC_16 port map( b(2) => B(3), b(1) => B(2), b(0) => B(1), A(31) =>
                           n205, A(30) => n205, A(29) => n205, A(28) => n205, 
                           A(27) => n205, A(26) => n205, A(25) => n205, A(24) 
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_34_port, p(31)
                           => q_0_1_33_port, p(30) => q_0_1_32_port, p(29) => 
                           q_0_1_31_port, p(28) => q_0_1_30_port, p(27) => 
                           q_0_1_29_port, p(26) => q_0_1_28_port, p(25) => 
                           q_0_1_27_port, p(24) => q_0_1_26_port, p(23) => 
                           q_0_1_25_port, p(22) => q_0_1_24_port, p(21) => 
                           q_0_1_23_port, p(20) => q_0_1_22_port, p(19) => 
                           q_0_1_21_port, p(18) => q_0_1_20_port, p(17) => 
                           q_0_1_19_port, p(16) => q_0_1_18_port, p(15) => 
                           q_0_1_17_port, p(14) => q_0_1_16_port, p(13) => 
                           q_0_1_15_port, p(12) => q_0_1_14_port, p(11) => 
                           q_0_1_13_port, p(10) => q_0_1_12_port, p(9) => 
                           q_0_1_11_port, p(8) => q_0_1_10_port, p(7) => 
                           q_0_1_9_port, p(6) => q_0_1_8_port, p(5) => 
                           q_0_1_7_port, p(4) => q_0_1_6_port, p(3) => 
                           q_0_1_5_port, p(2) => q_0_1_4_port, p(1) => 
                           q_0_1_3_port, p(0) => q_0_1_2_port);
   encI_3 : ENC_15 port map( b(2) => B(5), b(1) => B(4), b(0) => B(3), A(31) =>
                           n205, A(30) => n205, A(29) => n205, A(28) => n205, 
                           A(27) => n205, A(26) => n205, A(25) => n205, A(24) 
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_36_port, p(31)
                           => q_0_2_35_port, p(30) => q_0_2_34_port, p(29) => 
                           q_0_2_33_port, p(28) => q_0_2_32_port, p(27) => 
                           q_0_2_31_port, p(26) => q_0_2_30_port, p(25) => 
                           q_0_2_29_port, p(24) => q_0_2_28_port, p(23) => 
                           q_0_2_27_port, p(22) => q_0_2_26_port, p(21) => 
                           q_0_2_25_port, p(20) => q_0_2_24_port, p(19) => 
                           q_0_2_23_port, p(18) => q_0_2_22_port, p(17) => 
                           q_0_2_21_port, p(16) => q_0_2_20_port, p(15) => 
                           q_0_2_19_port, p(14) => q_0_2_18_port, p(13) => 
                           q_0_2_17_port, p(12) => q_0_2_16_port, p(11) => 
                           q_0_2_15_port, p(10) => q_0_2_14_port, p(9) => 
                           q_0_2_13_port, p(8) => q_0_2_12_port, p(7) => 
                           q_0_2_11_port, p(6) => q_0_2_10_port, p(5) => 
                           q_0_2_9_port, p(4) => q_0_2_8_port, p(3) => 
                           q_0_2_7_port, p(2) => q_0_2_6_port, p(1) => 
                           q_0_2_5_port, p(0) => q_0_2_4_port);
   encI_4 : ENC_14 port map( b(2) => B(7), b(1) => B(6), b(0) => B(5), A(31) =>
                           n205, A(30) => n205, A(29) => n205, A(28) => n205, 
                           A(27) => n205, A(26) => n205, A(25) => n205, A(24) 
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_38_port, p(31)
                           => q_0_1_37_port, p(30) => q_0_2_36_port, p(29) => 
                           q_0_3_35_port, p(28) => q_0_3_34_port, p(27) => 
                           q_0_3_33_port, p(26) => q_0_3_32_port, p(25) => 
                           q_0_3_31_port, p(24) => q_0_3_30_port, p(23) => 
                           q_0_3_29_port, p(22) => q_0_3_28_port, p(21) => 
                           q_0_3_27_port, p(20) => q_0_3_26_port, p(19) => 
                           q_0_3_25_port, p(18) => q_0_3_24_port, p(17) => 
                           q_0_3_23_port, p(16) => q_0_3_22_port, p(15) => 
                           q_0_3_21_port, p(14) => q_0_3_20_port, p(13) => 
                           q_0_3_19_port, p(12) => q_0_3_18_port, p(11) => 
                           q_0_3_17_port, p(10) => q_0_3_16_port, p(9) => 
                           q_0_3_15_port, p(8) => q_0_3_14_port, p(7) => 
                           q_0_3_13_port, p(6) => q_0_3_12_port, p(5) => 
                           q_0_3_11_port, p(4) => q_0_3_10_port, p(3) => 
                           q_0_3_9_port, p(2) => q_0_3_8_port, p(1) => 
                           q_0_3_7_port, p(0) => q_0_3_6_port);
   encI_5 : ENC_13 port map( b(2) => B(9), b(1) => B(8), b(0) => B(7), A(31) =>
                           n205, A(30) => n205, A(29) => n205, A(28) => n205, 
                           A(27) => n205, A(26) => n205, A(25) => n205, A(24) 
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_40_port, p(31)
                           => q_0_1_39_port, p(30) => q_0_2_38_port, p(29) => 
                           q_0_2_37_port, p(28) => q_0_3_36_port, p(27) => 
                           q_0_4_35_port, p(26) => q_0_4_34_port, p(25) => 
                           q_0_4_33_port, p(24) => q_0_4_32_port, p(23) => 
                           q_0_4_31_port, p(22) => q_0_4_30_port, p(21) => 
                           q_0_4_29_port, p(20) => q_0_4_28_port, p(19) => 
                           q_0_4_27_port, p(18) => q_0_4_26_port, p(17) => 
                           q_0_4_25_port, p(16) => q_0_4_24_port, p(15) => 
                           q_0_4_23_port, p(14) => q_0_4_22_port, p(13) => 
                           q_0_4_21_port, p(12) => q_0_4_20_port, p(11) => 
                           q_0_4_19_port, p(10) => q_0_4_18_port, p(9) => 
                           q_0_4_17_port, p(8) => q_0_4_16_port, p(7) => 
                           q_0_4_15_port, p(6) => q_0_4_14_port, p(5) => 
                           q_0_4_13_port, p(4) => q_0_4_12_port, p(3) => 
                           q_0_4_11_port, p(2) => q_0_4_10_port, p(1) => 
                           q_0_4_9_port, p(0) => q_0_4_8_port);
   encI_6 : ENC_12 port map( b(2) => B(11), b(1) => B(10), b(0) => B(9), A(31) 
                           => n205, A(30) => n205, A(29) => n205, A(28) => n205
                           , A(27) => n205, A(26) => n205, A(25) => n205, A(24)
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_42_port, p(31)
                           => q_0_1_41_port, p(30) => q_0_2_40_port, p(29) => 
                           q_0_2_39_port, p(28) => q_0_3_38_port, p(27) => 
                           q_0_3_37_port, p(26) => q_0_4_36_port, p(25) => 
                           q_0_5_35_port, p(24) => q_0_5_34_port, p(23) => 
                           q_0_5_33_port, p(22) => q_0_5_32_port, p(21) => 
                           q_0_5_31_port, p(20) => q_0_5_30_port, p(19) => 
                           q_0_5_29_port, p(18) => q_0_5_28_port, p(17) => 
                           q_0_5_27_port, p(16) => q_0_5_26_port, p(15) => 
                           q_0_5_25_port, p(14) => q_0_5_24_port, p(13) => 
                           q_0_5_23_port, p(12) => q_0_5_22_port, p(11) => 
                           q_0_5_21_port, p(10) => q_0_5_20_port, p(9) => 
                           q_0_5_19_port, p(8) => q_0_5_18_port, p(7) => 
                           q_0_5_17_port, p(6) => q_0_5_16_port, p(5) => 
                           q_0_5_15_port, p(4) => q_0_5_14_port, p(3) => 
                           q_0_5_13_port, p(2) => q_0_5_12_port, p(1) => 
                           q_0_5_11_port, p(0) => q_0_5_10_port);
   encI_7 : ENC_11 port map( b(2) => B(13), b(1) => B(12), b(0) => B(11), A(31)
                           => n205, A(30) => n205, A(29) => n205, A(28) => n205
                           , A(27) => n205, A(26) => n205, A(25) => n205, A(24)
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_44_port, p(31)
                           => q_0_1_43_port, p(30) => q_0_2_42_port, p(29) => 
                           q_0_2_41_port, p(28) => q_0_3_40_port, p(27) => 
                           q_0_3_39_port, p(26) => q_0_4_38_port, p(25) => 
                           q_0_4_37_port, p(24) => q_0_5_36_port, p(23) => 
                           q_0_6_35_port, p(22) => q_0_6_34_port, p(21) => 
                           q_0_6_33_port, p(20) => q_0_6_32_port, p(19) => 
                           q_0_6_31_port, p(18) => q_0_6_30_port, p(17) => 
                           q_0_6_29_port, p(16) => q_0_6_28_port, p(15) => 
                           q_0_6_27_port, p(14) => q_0_6_26_port, p(13) => 
                           q_0_6_25_port, p(12) => q_0_6_24_port, p(11) => 
                           q_0_6_23_port, p(10) => q_0_6_22_port, p(9) => 
                           q_0_6_21_port, p(8) => q_0_6_20_port, p(7) => 
                           q_0_6_19_port, p(6) => q_0_6_18_port, p(5) => 
                           q_0_6_17_port, p(4) => q_0_6_16_port, p(3) => 
                           q_0_6_15_port, p(2) => q_0_6_14_port, p(1) => 
                           q_0_6_13_port, p(0) => q_0_6_12_port);
   encI_8 : ENC_10 port map( b(2) => B(15), b(1) => B(14), b(0) => B(13), A(31)
                           => n205, A(30) => n205, A(29) => n205, A(28) => n205
                           , A(27) => n205, A(26) => n205, A(25) => n205, A(24)
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_46_port, p(31)
                           => q_0_1_45_port, p(30) => q_0_2_44_port, p(29) => 
                           q_0_2_43_port, p(28) => q_0_3_42_port, p(27) => 
                           q_0_3_41_port, p(26) => q_0_4_40_port, p(25) => 
                           q_0_4_39_port, p(24) => q_0_5_38_port, p(23) => 
                           q_0_5_37_port, p(22) => q_0_6_36_port, p(21) => 
                           q_0_7_35_port, p(20) => q_0_7_34_port, p(19) => 
                           q_0_7_33_port, p(18) => q_0_7_32_port, p(17) => 
                           q_0_7_31_port, p(16) => q_0_7_30_port, p(15) => 
                           q_0_7_29_port, p(14) => q_0_7_28_port, p(13) => 
                           q_0_7_27_port, p(12) => q_0_7_26_port, p(11) => 
                           q_0_7_25_port, p(10) => q_0_7_24_port, p(9) => 
                           q_0_7_23_port, p(8) => q_0_7_22_port, p(7) => 
                           q_0_7_21_port, p(6) => q_0_7_20_port, p(5) => 
                           q_0_7_19_port, p(4) => q_0_7_18_port, p(3) => 
                           q_0_7_17_port, p(2) => q_0_7_16_port, p(1) => 
                           q_0_7_15_port, p(0) => q_0_7_14_port);
   encI_9 : ENC_9 port map( b(2) => B(17), b(1) => B(16), b(0) => B(15), A(31) 
                           => n205, A(30) => n205, A(29) => n205, A(28) => n205
                           , A(27) => n205, A(26) => n205, A(25) => n205, A(24)
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2251, p(31) => 
                           q_0_1_47_port, p(30) => q_0_2_46_port, p(29) => 
                           q_0_2_45_port, p(28) => q_0_3_44_port, p(27) => 
                           q_0_3_43_port, p(26) => q_0_4_42_port, p(25) => 
                           q_0_4_41_port, p(24) => q_0_5_40_port, p(23) => 
                           q_0_5_39_port, p(22) => q_0_6_38_port, p(21) => 
                           q_0_6_37_port, p(20) => q_0_7_36_port, p(19) => 
                           q_0_8_35_port, p(18) => q_0_8_34_port, p(17) => 
                           q_0_8_33_port, p(16) => q_0_8_32_port, p(15) => 
                           q_0_8_31_port, p(14) => q_0_8_30_port, p(13) => 
                           q_0_8_29_port, p(12) => q_0_8_28_port, p(11) => 
                           q_0_8_27_port, p(10) => q_0_8_26_port, p(9) => 
                           q_0_8_25_port, p(8) => q_0_8_24_port, p(7) => 
                           q_0_8_23_port, p(6) => q_0_8_22_port, p(5) => 
                           q_0_8_21_port, p(4) => q_0_8_20_port, p(3) => 
                           q_0_8_19_port, p(2) => q_0_8_18_port, p(1) => 
                           q_0_8_17_port, p(0) => q_0_8_16_port);
   encI_10 : ENC_8 port map( b(2) => B(19), b(1) => B(18), b(0) => B(17), A(31)
                           => n205, A(30) => n205, A(29) => n205, A(28) => n205
                           , A(27) => n205, A(26) => n205, A(25) => n205, A(24)
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2252, p(31) => 
                           n_2253, p(30) => n_2254, p(29) => q_0_2_47_port, 
                           p(28) => q_0_3_46_port, p(27) => q_0_3_45_port, 
                           p(26) => q_0_4_44_port, p(25) => q_0_4_43_port, 
                           p(24) => q_0_5_42_port, p(23) => q_0_5_41_port, 
                           p(22) => q_0_6_40_port, p(21) => q_0_6_39_port, 
                           p(20) => q_0_7_38_port, p(19) => q_0_7_37_port, 
                           p(18) => q_0_8_36_port, p(17) => q_0_9_35_port, 
                           p(16) => q_0_9_34_port, p(15) => q_0_9_33_port, 
                           p(14) => q_0_9_32_port, p(13) => q_0_9_31_port, 
                           p(12) => q_0_9_30_port, p(11) => q_0_9_29_port, 
                           p(10) => q_0_9_28_port, p(9) => q_0_9_27_port, p(8) 
                           => q_0_9_26_port, p(7) => q_0_9_25_port, p(6) => 
                           q_0_9_24_port, p(5) => q_0_9_23_port, p(4) => 
                           q_0_9_22_port, p(3) => q_0_9_21_port, p(2) => 
                           q_0_9_20_port, p(1) => q_0_9_19_port, p(0) => 
                           q_0_9_18_port);
   encI_11 : ENC_7 port map( b(2) => B(21), b(1) => B(20), b(0) => B(19), A(31)
                           => n205, A(30) => n205, A(29) => n205, A(28) => n205
                           , A(27) => n205, A(26) => n205, A(25) => n205, A(24)
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2255, p(31) => 
                           n_2256, p(30) => n_2257, p(29) => n_2258, p(28) => 
                           n_2259, p(27) => q_0_3_47_port, p(26) => 
                           q_0_4_46_port, p(25) => q_0_4_45_port, p(24) => 
                           q_0_5_44_port, p(23) => q_0_5_43_port, p(22) => 
                           q_0_6_42_port, p(21) => q_0_6_41_port, p(20) => 
                           q_0_7_40_port, p(19) => q_0_7_39_port, p(18) => 
                           q_0_8_38_port, p(17) => q_0_8_37_port, p(16) => 
                           q_0_9_36_port, p(15) => q_0_10_35_port, p(14) => 
                           q_0_10_34_port, p(13) => q_0_10_33_port, p(12) => 
                           q_0_10_32_port, p(11) => q_0_10_31_port, p(10) => 
                           q_0_10_30_port, p(9) => q_0_10_29_port, p(8) => 
                           q_0_10_28_port, p(7) => q_0_10_27_port, p(6) => 
                           q_0_10_26_port, p(5) => q_0_10_25_port, p(4) => 
                           q_0_10_24_port, p(3) => q_0_10_23_port, p(2) => 
                           q_0_10_22_port, p(1) => q_0_10_21_port, p(0) => 
                           q_0_10_20_port);
   encI_12 : ENC_6 port map( b(2) => B(23), b(1) => B(22), b(0) => B(21), A(31)
                           => n205, A(30) => n205, A(29) => n205, A(28) => n205
                           , A(27) => n205, A(26) => n205, A(25) => n205, A(24)
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2260, p(31) => 
                           n_2261, p(30) => n_2262, p(29) => n_2263, p(28) => 
                           n_2264, p(27) => n_2265, p(26) => n_2266, p(25) => 
                           q_0_4_47_port, p(24) => q_0_5_46_port, p(23) => 
                           q_0_5_45_port, p(22) => q_0_6_44_port, p(21) => 
                           q_0_6_43_port, p(20) => q_0_7_42_port, p(19) => 
                           q_0_7_41_port, p(18) => q_0_8_40_port, p(17) => n191
                           , p(16) => q_0_9_38_port, p(15) => q_0_9_37_port, 
                           p(14) => q_0_10_36_port, p(13) => q_0_11_35_port, 
                           p(12) => q_0_11_34_port, p(11) => q_0_11_33_port, 
                           p(10) => q_0_11_32_port, p(9) => q_0_11_31_port, 
                           p(8) => q_0_11_30_port, p(7) => q_0_11_29_port, p(6)
                           => q_0_11_28_port, p(5) => q_0_11_27_port, p(4) => 
                           q_0_11_26_port, p(3) => q_0_11_25_port, p(2) => 
                           q_0_11_24_port, p(1) => q_0_11_23_port, p(0) => 
                           q_0_11_22_port);
   encI_13 : ENC_5 port map( b(2) => n213, b(1) => n214, b(0) => B(23), A(31) 
                           => n205, A(30) => n205, A(29) => n205, A(28) => n205
                           , A(27) => n205, A(26) => n205, A(25) => n205, A(24)
                           => n205, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2267, p(31) => 
                           n_2268, p(30) => n_2269, p(29) => n_2270, p(28) => 
                           n_2271, p(27) => n_2272, p(26) => n_2273, p(25) => 
                           n_2274, p(24) => n_2275, p(23) => q_0_5_47_port, 
                           p(22) => q_0_6_46_port, p(21) => q_0_6_45_port, 
                           p(20) => q_0_7_44_port, p(19) => q_0_7_43_port, 
                           p(18) => q_0_8_42_port, p(17) => q_0_8_41_port, 
                           p(16) => q_0_9_40_port, p(15) => q_0_9_39_port, 
                           p(14) => q_0_10_38_port, p(13) => q_0_10_37_port, 
                           p(12) => q_0_11_36_port, p(11) => q_0_12_35_port, 
                           p(10) => q_0_12_34_port, p(9) => q_0_12_33_port, 
                           p(8) => q_0_12_32_port, p(7) => q_0_12_31_port, p(6)
                           => q_0_12_30_port, p(5) => q_0_12_29_port, p(4) => 
                           q_0_12_28_port, p(3) => q_0_12_27_port, p(2) => 
                           q_0_12_26_port, p(1) => q_0_12_25_port, p(0) => 
                           q_0_12_24_port);
   encI_14 : ENC_4 port map( b(2) => n211, b(1) => n212, b(0) => n213, A(31) =>
                           n205, A(30) => n205, A(29) => n205, A(28) => n205, 
                           A(27) => n205, A(26) => n205, A(25) => n205, A(24) 
                           => n205, A(23) => n120, A(22) => n121, A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           net102814, A(14) => net102815, A(13) => net102816, 
                           A(12) => net102817, A(11) => net102818, A(10) => 
                           net102819, A(9) => net102820, A(8) => net102821, 
                           A(7) => net102822, A(6) => net102823, A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), clk => clk, p_32_port => n_2276,
                           p_31_port => n_2277, p_30_port => n_2278, p_29_port 
                           => n_2279, p_28_port => n_2280, p_27_port => n_2281,
                           p_26_port => n_2282, p_25_port => n_2283, p_24_port 
                           => n_2284, p_23_port => n_2285, p_22_port => n_2286,
                           p_21_port => q_0_6_47_port, p_20_port => 
                           q_0_7_46_port, p_19_port => q_0_7_45_port, p_18_port
                           => q_0_8_44_port, p_17_port => q_0_8_43_port, 
                           p_15_port => n_2287, p_14_port => n_2288, p_13_port 
                           => n_2289, p_12_port => n_2290, p_11_port => n_2291,
                           p_10_port => n_2292, p_9_port => n_2293, p_8_port =>
                           n_2294, p_7_port => n_2295, p_6_BAR => 
                           q_0_13_32_port, p_5_port => q_0_13_31_port, p_4_port
                           => q_0_13_30_port, p_3_port => q_0_13_29_port, 
                           p_2_port => q_0_13_28_port, p_1_port => 
                           q_0_13_27_port, p_0_port => q_0_13_26_port, p_16_BAR
                           => q_0_9_42_port);
   encI_15 : ENC_3 port map( b(2) => n209, b(1) => n210, b(0) => n211, A(31) =>
                           n205, A(30) => n205, A(29) => n205, A(28) => n205, 
                           A(27) => n205, A(26) => n205, A(25) => n205, A(24) 
                           => n205, A(23) => n122, A(22) => n123, A(21) => n124
                           , A(20) => n125, A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => net102802, 
                           A(14) => net102803, A(13) => net102804, A(12) => 
                           net102805, A(11) => net102806, A(10) => net102807, 
                           A(9) => net102808, A(8) => net102809, A(7) => 
                           net102810, A(6) => net102811, A(5) => net102812, 
                           A(4) => net102813, A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), clk => clk, p_32_port => 
                           n_2296, p_31_port => n_2297, p_30_port => n_2298, 
                           p_29_port => n_2299, p_28_port => n_2300, p_27_port 
                           => n_2301, p_26_port => n_2302, p_25_port => n_2303,
                           p_24_port => n_2304, p_23_port => n_2305, p_22_port 
                           => n_2306, p_21_port => n_2307, p_20_port => n_2308,
                           p_19_port => q_0_7_47_port, p_18_port => 
                           q_0_8_46_port, p_17_port => q_0_8_45_port, p_15_port
                           => n_2309, p_14_port => n_2310, p_13_port => n_2311,
                           p_12_port => n_2312, p_11_port => n_2313, p_10_port 
                           => n_2314, p_9_port => n_2315, p_8_port => n_2316, 
                           p_7_port => n_2317, p_6_port => n_2318, p_5_port => 
                           n_2319, p_4_BAR => q_0_14_32_port, p_3_port => 
                           q_0_14_31_port, p_2_port => q_0_14_30_port, p_1_port
                           => q_0_14_29_port, p_0_port => q_0_14_28_port, 
                           p_16_BAR => q_0_9_44_port);
   encI_16 : ENC_2 port map( b(2) => n207, b(1) => n208, b(0) => n209, A(31) =>
                           n205, A(30) => n205, A(29) => n205, A(28) => n205, 
                           A(27) => n205, A(26) => n205, A(25) => n205, A(24) 
                           => n205, A(23) => n126, A(22) => n127, A(21) => n128
                           , A(20) => n129, A(19) => n130, A(18) => n131, A(17)
                           => A(17), A(16) => A(16), A(15) => net102786, A(14) 
                           => net102787, A(13) => net102788, A(12) => net102789
                           , A(11) => net102790, A(10) => net102791, A(9) => 
                           net102792, A(8) => net102793, A(7) => net102794, 
                           A(6) => net102795, A(5) => net102796, A(4) => 
                           net102797, A(3) => net102798, A(2) => net102799, 
                           A(1) => net102800, A(0) => net102801, clk => clk, 
                           p_32_port => n_2320, p_31_port => n_2321, p_30_port 
                           => n_2322, p_29_port => n_2323, p_28_port => n_2324,
                           p_27_port => n_2325, p_26_port => n_2326, p_25_port 
                           => n_2327, p_24_port => n_2328, p_23_port => n_2329,
                           p_22_port => n_2330, p_21_port => n_2331, p_20_port 
                           => n_2332, p_19_port => n_2333, p_18_port => n_2334,
                           p_17_port => q_0_8_47_port, p_16_BAR => 
                           q_0_9_46_port, p_15_port => n_2335, p_14_port => 
                           n_2336, p_13_port => n_2337, p_12_port => n_2338, 
                           p_11_port => n_2339, p_10_port => n_2340, p_9_port 
                           => n_2341, p_8_port => n_2342, p_7_port => n_2343, 
                           p_6_port => n_2344, p_5_port => n_2345, p_4_port => 
                           n_2346, p_3_port => n_2347, p_2_port => n_2348, 
                           p_1_port => n_2349, p_0_port => n_2350);
   encI_17 : ENC_1 port map( b(2) => X_Logic0_port, b(1) => X_Logic0_port, b(0)
                           => n207, A(31) => n205, A(30) => n205, A(29) => n205
                           , A(28) => n205, A(27) => n205, A(26) => n205, A(25)
                           => n205, A(24) => n205, A(23) => n132, A(22) => n133
                           , A(21) => n134, A(20) => n135, A(19) => n136, A(18)
                           => n137, A(17) => n138, A(16) => n139, A(15) => 
                           A(15), A(14) => A(14), A(13) => net102772, A(12) => 
                           net102773, A(11) => net102774, A(10) => net102775, 
                           A(9) => net102776, A(8) => net102777, A(7) => 
                           net102778, A(6) => net102779, A(5) => net102780, 
                           A(4) => net102781, A(3) => net102782, A(2) => 
                           net102783, A(1) => net102784, A(0) => net102785, clk
                           => clk, p_32_port => n_2351, p_31_port => n_2352, 
                           p_30_port => n_2353, p_29_port => n_2354, p_28_port 
                           => n_2355, p_27_port => n_2356, p_26_port => n_2357,
                           p_25_port => n_2358, p_24_port => n_2359, p_23_port 
                           => n_2360, p_22_port => n_2361, p_21_port => n_2362,
                           p_20_port => n_2363, p_19_port => n_2364, p_18_port 
                           => n_2365, p_17_port => n_2366, p_16_port => n_2367,
                           p_15_port => q_0_9_47_port, p_14_BAR => 
                           q_0_10_46_port, p_13_port => n_2368, p_12_port => 
                           n_2369, p_11_port => n_2370, p_10_port => n_2371, 
                           p_9_port => n_2372, p_8_port => n_2373, p_7_port => 
                           n_2374, p_6_port => n_2375, p_5_port => n_2376, 
                           p_4_port => n_2377, p_3_port => n_2378, p_2_port => 
                           n_2379, p_1_port => n_2380, p_0_port => n_2381);
   HA_R_0_0_24 : HA_0 port map( A => q_0_0_24_port, B => q_0_1_24_port, S => 
                           q_1_0_24_port, C => q_1_1_25_port);
   HA_R_0_0_25 : HA_43 port map( A => q_0_0_25_port, B => q_0_1_25_port, S => 
                           q_1_0_25_port, C => q_1_1_26_port);
   FA_C_0_0_26 : FA_0 port map( A => q_0_0_26_port, B => q_0_1_26_port, Ci => 
                           q_0_2_26_port, S => q_1_0_26_port, Co => 
                           q_1_1_27_port);
   FA_C_0_0_27 : FA_607 port map( A => q_0_0_27_port, B => q_0_1_27_port, Ci =>
                           q_0_2_27_port, S => q_1_0_27_port, Co => 
                           q_1_1_28_port);
   FA_C_0_0_28 : FA_606 port map( A => q_0_0_28_port, B => q_0_1_28_port, Ci =>
                           q_0_2_28_port, S => q_1_0_28_port, Co => 
                           q_1_1_29_port);
   FA_C_0_0_29 : FA_605 port map( A => q_0_0_29_port, B => q_0_1_29_port, Ci =>
                           q_0_2_29_port, S => q_1_0_29_port, Co => 
                           q_1_1_30_port);
   FA_C_0_0_30 : FA_604 port map( A => q_0_0_30_port, B => q_0_1_30_port, Ci =>
                           q_0_2_30_port, S => q_1_0_30_port, Co => 
                           q_1_1_31_port);
   FA_C_0_0_31 : FA_603 port map( A => q_0_0_31_port, B => q_0_1_31_port, Ci =>
                           q_0_2_31_port, S => q_1_0_31_port, Co => 
                           q_1_1_32_port);
   FA_C_0_0_32 : FA_602 port map( A => q_0_0_32_port, B => q_0_1_32_port, Ci =>
                           q_0_2_32_port, S => q_1_0_32_port, Co => 
                           q_1_1_33_port);
   FA_C_0_0_33 : FA_601 port map( A => B(1), B => q_0_1_33_port, Ci => 
                           q_0_2_33_port, S => q_1_0_33_port, Co => 
                           q_1_1_34_port);
   FA_C_0_0_34 : FA_600 port map( B => q_0_1_34_port, Ci => q_0_2_34_port, S =>
                           q_1_0_34_port, Co => q_1_1_35_port, A_BAR => n95);
   FA_C_0_0_35 : FA_599 port map( A => n95, Ci => q_0_2_35_port, S => 
                           q_1_0_35_port, Co => q_1_1_36_port, B_BAR => B(3));
   FA_C_0_0_36 : FA_598 port map( A => X_Logic1_port, B => q_0_1_36_port, Ci =>
                           q_0_2_36_port, S => q_1_0_36_port, Co => 
                           q_1_1_37_port);
   FA_C_0_0_37 : FA_597 port map( A => n93, B => q_0_1_37_port, Ci => 
                           q_0_2_37_port, S => q_1_0_37_port, Co => 
                           q_1_1_38_port);
   FA_C_0_0_38 : FA_596 port map( A => X_Logic1_port, B => q_0_1_38_port, Ci =>
                           q_0_2_38_port, S => q_1_0_38_port, Co => 
                           q_1_1_39_port);
   FA_C_0_0_39 : FA_595 port map( A => n92, B => q_0_1_39_port, Ci => 
                           q_0_2_39_port, S => q_1_0_39_port, Co => 
                           q_1_1_40_port);
   FA_C_0_0_40 : FA_594 port map( A => X_Logic1_port, B => q_0_1_40_port, Ci =>
                           q_0_2_40_port, S => q_1_0_40_port, Co => 
                           q_1_1_41_port);
   FA_C_0_0_41 : FA_593 port map( A => n91, B => q_0_1_41_port, Ci => 
                           q_0_2_41_port, S => q_1_0_41_port, Co => 
                           q_1_1_42_port);
   HA_L_0_0_42 : HA_42 port map( A => X_Logic1_port, B => q_0_1_42_port, S => 
                           q_1_0_42_port, C => q_1_0_43_port);
   HA_R_0_3_26 : HA_41 port map( A => q_0_3_26_port, B => q_0_4_26_port, S => 
                           q_1_2_26_port, C => q_1_3_27_port);
   HA_R_0_3_27 : HA_40 port map( A => q_0_3_27_port, B => q_0_4_27_port, S => 
                           q_1_2_27_port, C => q_1_3_28_port);
   FA_C_0_3_28 : FA_592 port map( A => q_0_3_28_port, B => q_0_4_28_port, Ci =>
                           q_0_5_28_port, S => q_1_2_28_port, Co => 
                           q_1_3_29_port);
   FA_C_0_3_29 : FA_591 port map( A => q_0_3_29_port, B => q_0_4_29_port, Ci =>
                           q_0_5_29_port, S => q_1_2_29_port, Co => n190);
   FA_C_0_3_30 : FA_590 port map( A => q_0_3_30_port, B => q_0_4_30_port, Ci =>
                           q_0_5_30_port, S => q_1_2_30_port, Co => 
                           q_1_3_31_port);
   FA_C_0_3_31 : FA_589 port map( A => q_0_3_31_port, B => q_0_4_31_port, Ci =>
                           q_0_5_31_port, S => n182, Co => q_1_3_32_port);
   FA_C_0_3_32 : FA_588 port map( A => q_0_3_32_port, B => q_0_4_32_port, Ci =>
                           q_0_5_32_port, S => q_1_2_32_port, Co => 
                           q_1_3_33_port);
   FA_C_0_3_33 : FA_587 port map( A => q_0_3_33_port, B => q_0_4_33_port, Ci =>
                           q_0_5_33_port, S => q_1_2_33_port, Co => 
                           q_1_3_34_port);
   FA_C_0_3_34 : FA_586 port map( A => q_0_3_34_port, B => q_0_4_34_port, Ci =>
                           q_0_5_34_port, S => q_1_2_34_port, Co => 
                           q_1_3_35_port);
   FA_C_0_3_35 : FA_585 port map( A => q_0_3_35_port, B => q_0_4_35_port, Ci =>
                           q_0_5_35_port, S => q_1_2_35_port, Co => 
                           q_1_3_36_port);
   FA_C_0_3_36 : FA_584 port map( A => q_0_3_36_port, B => q_0_4_36_port, Ci =>
                           q_0_5_36_port, S => n181, Co => q_1_3_37_port);
   FA_C_0_3_37 : FA_583 port map( A => q_0_3_37_port, B => q_0_4_37_port, Ci =>
                           q_0_5_37_port, S => q_1_2_37_port, Co => 
                           q_1_3_38_port);
   FA_C_0_3_38 : FA_582 port map( A => q_0_3_38_port, B => q_0_4_38_port, Ci =>
                           q_0_5_38_port, S => q_1_2_38_port, Co => 
                           q_1_3_39_port);
   FA_C_0_3_39 : FA_581 port map( A => q_0_3_39_port, B => q_0_4_39_port, Ci =>
                           q_0_5_39_port, S => q_1_2_39_port, Co => 
                           q_1_3_40_port);
   HA_L_0_3_40 : HA_39 port map( A => q_0_3_40_port, B => q_0_4_40_port, S => 
                           q_1_2_40_port, C => q_1_2_41_port);
   HA_R_0_6_28 : HA_38 port map( A => q_0_6_28_port, B => q_0_7_28_port, S => 
                           q_1_4_28_port, C => q_1_5_29_port);
   HA_R_0_6_29 : HA_37 port map( A => q_0_6_29_port, B => q_0_7_29_port, S => 
                           q_1_4_29_port, C => q_1_5_30_port);
   FA_C_0_6_30 : FA_580 port map( A => q_0_6_30_port, B => q_0_7_30_port, Ci =>
                           q_0_8_30_port, S => q_1_4_30_port, Co => 
                           q_1_5_31_port);
   FA_C_0_6_31 : FA_579 port map( A => q_0_6_31_port, B => q_0_7_31_port, Ci =>
                           q_0_8_31_port, S => q_1_4_31_port, Co => 
                           q_1_5_32_port);
   FA_C_0_6_32 : FA_578 port map( A => q_0_6_32_port, B => q_0_7_32_port, Ci =>
                           q_0_8_32_port, S => q_1_4_32_port, Co => 
                           q_1_5_33_port);
   FA_C_0_6_33 : FA_577 port map( A => q_0_6_33_port, B => q_0_7_33_port, Ci =>
                           q_0_8_33_port, S => q_1_4_33_port, Co => 
                           q_1_5_34_port);
   FA_C_0_6_34 : FA_576 port map( A => q_0_6_34_port, B => q_0_7_34_port, Ci =>
                           q_0_8_34_port, S => q_1_4_34_port, Co => n184);
   FA_C_0_6_35 : FA_575 port map( A => q_0_6_35_port, B => q_0_7_35_port, Ci =>
                           q_0_8_35_port, S => q_1_4_35_port, Co => 
                           q_1_5_36_port);
   FA_C_0_6_36 : FA_574 port map( A => q_0_6_36_port, B => q_0_7_36_port, Ci =>
                           q_0_8_36_port, S => q_1_4_36_port, Co => 
                           q_1_5_37_port);
   FA_C_0_6_37 : FA_573 port map( A => q_0_6_37_port, B => q_0_7_37_port, Ci =>
                           q_0_8_37_port, S => q_1_4_37_port, Co => 
                           q_1_5_38_port);
   HA_L_0_6_38 : HA_36 port map( A => q_0_6_38_port, B => q_0_7_38_port, S => 
                           q_1_4_38_port, C => q_1_4_39_port);
   HA_R_0_9_30 : HA_35 port map( A => q_0_9_30_port, B => q_0_10_30_port, S => 
                           n189, C => q_1_7_31_port);
   HA_R_0_9_31 : HA_34 port map( A => q_0_9_31_port, B => q_0_10_31_port, S => 
                           q_1_6_31_port, C => q_1_7_32_port);
   FA_C_0_9_32 : FA_572 port map( A => q_0_9_32_port, B => q_0_10_32_port, Ci 
                           => q_0_11_32_port, S => q_1_6_32_port, Co => 
                           q_1_7_33_port);
   FA_C_0_9_33 : FA_571 port map( A => q_0_9_33_port, B => q_0_10_33_port, Ci 
                           => q_0_11_33_port, S => q_1_6_33_port, Co => 
                           q_1_7_34_port);
   FA_C_0_9_34 : FA_570 port map( A => q_0_9_34_port, B => q_0_10_34_port, Ci 
                           => q_0_11_34_port, S => q_1_6_34_port, Co => 
                           q_1_7_35_port);
   FA_C_0_9_35 : FA_569 port map( A => q_0_9_35_port, B => q_0_10_35_port, Ci 
                           => q_0_11_35_port, S => q_1_6_35_port, Co => n179);
   HA_L_0_9_36 : HA_33 port map( A => q_0_9_36_port, B => q_0_10_36_port, S => 
                           q_1_6_36_port, C => q_1_6_37_port);
   HA_R_1_0_16 : HA_32 port map( A => q_0_0_16_port, B => q_0_1_16_port, S => 
                           q_2_0_16_port, C => q_2_1_17_port);
   HA_R_1_0_17 : HA_31 port map( A => q_0_0_17_port, B => q_0_1_17_port, S => 
                           q_2_0_17_port, C => q_2_1_18_port);
   FA_C_1_0_18 : FA_568 port map( A => q_0_0_18_port, B => q_0_1_18_port, Ci =>
                           q_0_2_18_port, S => q_2_0_18_port, Co => 
                           q_2_1_19_port);
   FA_C_1_0_19 : FA_567 port map( A => q_0_0_19_port, B => q_0_1_19_port, Ci =>
                           q_0_2_19_port, S => q_2_0_19_port, Co => 
                           q_2_1_20_port);
   FA_C_1_0_20 : FA_566 port map( A => q_0_0_20_port, B => q_0_1_20_port, Ci =>
                           q_0_2_20_port, S => q_2_0_20_port, Co => 
                           q_2_1_21_port);
   FA_C_1_0_21 : FA_565 port map( A => q_0_0_21_port, B => q_0_1_21_port, Ci =>
                           q_0_2_21_port, S => q_2_0_21_port, Co => 
                           q_2_1_22_port);
   FA_C_1_0_22 : FA_564 port map( A => q_0_0_22_port, B => q_0_1_22_port, Ci =>
                           q_0_2_22_port, S => q_2_0_22_port, Co => 
                           q_2_1_23_port);
   FA_C_1_0_23 : FA_563 port map( A => q_0_0_23_port, B => q_0_1_23_port, Ci =>
                           q_0_2_23_port, S => q_2_0_23_port, Co => 
                           q_2_1_24_port);
   FA_C_1_0_24 : FA_562 port map( A => q_1_0_24_port, B => q_0_2_24_port, Ci =>
                           q_0_3_24_port, S => q_2_0_24_port, Co => 
                           q_2_1_25_port);
   FA_C_1_0_25 : FA_561 port map( A => q_1_0_25_port, B => q_1_1_25_port, Ci =>
                           q_0_2_25_port, S => q_2_0_25_port, Co => 
                           q_2_1_26_port);
   FA_C_1_0_26 : FA_560 port map( A => q_1_0_26_port, B => q_1_1_26_port, Ci =>
                           q_1_2_26_port, S => q_2_0_26_port, Co => 
                           q_2_1_27_port);
   FA_C_1_0_27 : FA_559 port map( A => q_1_0_27_port, B => q_1_1_27_port, Ci =>
                           q_1_2_27_port, S => q_2_0_27_port, Co => 
                           q_2_1_28_port);
   FA_C_1_0_28 : FA_558 port map( A => q_1_0_28_port, B => q_1_1_28_port, Ci =>
                           q_1_2_28_port, S => q_2_0_28_port, Co => 
                           q_2_1_29_port);
   FA_C_1_0_29 : FA_557 port map( A => q_1_0_29_port, B => q_1_1_29_port, Ci =>
                           q_1_2_29_port, S => q_2_0_29_port, Co => 
                           q_2_1_30_port);
   FA_C_1_0_30 : FA_556 port map( A => q_1_0_30_port, B => q_1_1_30_port, Ci =>
                           q_1_2_30_port, S => q_2_0_30_port, Co => 
                           q_2_1_31_port);
   FA_C_1_0_31 : FA_555 port map( A => q_1_0_31_port, B => q_1_1_31_port, Ci =>
                           n182, S => q_2_0_31_port, Co => q_2_1_32_port);
   FA_C_1_0_32 : FA_554 port map( A => q_1_0_32_port, B => q_1_1_32_port, Ci =>
                           q_1_2_32_port, S => q_2_0_32_port, Co => 
                           q_2_1_33_port);
   FA_C_1_0_33 : FA_553 port map( A => q_1_0_33_port, B => q_1_1_33_port, Ci =>
                           q_1_2_33_port, S => q_2_0_33_port, Co => 
                           q_2_1_34_port);
   FA_C_1_0_34 : FA_552 port map( A => q_1_0_34_port, B => q_1_1_34_port, Ci =>
                           q_1_2_34_port, S => q_2_0_34_port, Co => 
                           q_2_1_35_port, clk => clk);
   FA_C_1_0_35 : FA_551 port map( A => q_1_0_35_port, B => q_1_1_35_port, Ci =>
                           q_1_2_35_port, S => q_2_0_35_port, Co => 
                           q_2_1_36_port);
   FA_C_1_0_36 : FA_550 port map( A => q_1_0_36_port, B => q_1_1_36_port, Ci =>
                           n181, S => q_2_0_36_port, Co => q_2_1_37_port);
   FA_C_1_0_37 : FA_549 port map( A => q_1_0_37_port, B => q_1_1_37_port, Ci =>
                           q_1_2_37_port, S => q_2_0_37_port, Co => 
                           q_2_1_38_port);
   FA_C_1_0_38 : FA_548 port map( A => q_1_0_38_port, B => q_1_1_38_port, Ci =>
                           q_1_2_38_port, S => q_2_0_38_port, Co => 
                           q_2_1_39_port);
   FA_C_1_0_39 : FA_547 port map( A => q_1_0_39_port, B => q_1_1_39_port, Ci =>
                           q_1_2_39_port, S => q_2_0_39_port, Co => 
                           q_2_1_40_port);
   FA_C_1_0_40 : FA_546 port map( A => q_1_0_40_port, B => q_1_1_40_port, Ci =>
                           q_1_2_40_port, S => q_2_0_40_port, Co => 
                           q_2_1_41_port);
   FA_C_1_0_41 : FA_545 port map( A => q_1_0_41_port, B => q_1_1_41_port, Ci =>
                           q_1_2_41_port, S => q_2_0_41_port, Co => 
                           q_2_1_42_port);
   FA_C_1_0_42 : FA_544 port map( A => q_1_0_42_port, B => q_1_1_42_port, Ci =>
                           q_0_2_42_port, S => q_2_0_42_port, Co => 
                           q_2_1_43_port);
   FA_C_1_0_43 : FA_543 port map( A => q_1_0_43_port, Ci => q_0_1_43_port, S =>
                           q_2_0_43_port, Co => q_2_1_44_port, B_BAR => B(11));
   FA_C_1_0_44 : FA_542 port map( A => X_Logic1_port, B => q_0_1_44_port, Ci =>
                           q_0_2_44_port, S => q_2_0_44_port, Co => 
                           q_2_1_45_port);
   FA_C_1_0_45 : FA_541 port map( B => q_0_1_45_port, Ci => q_0_2_45_port, S =>
                           q_2_0_45_port, Co => q_2_1_46_port, A_BAR => B(13));
   FA_C_1_0_46 : FA_540 port map( A => X_Logic1_port, B => q_0_1_46_port, Ci =>
                           q_0_2_46_port, S => q_2_0_46_port, Co => 
                           q_2_1_47_port);
   FA_C_1_0_47 : FA_539 port map( B => q_0_1_47_port, Ci => q_0_2_47_port, S =>
                           q_2_0_47_port, Co => n_2382, A_BAR => B(15));
   HA_R_1_3_18 : HA_29 port map( A => q_0_3_18_port, B => q_0_4_18_port, S => 
                           q_2_2_18_port, C => q_2_3_19_port);
   HA_R_1_3_19 : HA_28 port map( A => q_0_3_19_port, B => q_0_4_19_port, S => 
                           q_2_2_19_port, C => q_2_3_20_port);
   FA_C_1_3_20 : FA_536 port map( A => q_0_3_20_port, B => q_0_4_20_port, Ci =>
                           q_0_5_20_port, S => q_2_2_20_port, Co => 
                           q_2_3_21_port);
   FA_C_1_3_21 : FA_535 port map( A => q_0_3_21_port, B => q_0_4_21_port, Ci =>
                           q_0_5_21_port, S => q_2_2_21_port, Co => 
                           q_2_3_22_port);
   FA_C_1_3_22 : FA_534 port map( A => q_0_3_22_port, B => q_0_4_22_port, Ci =>
                           q_0_5_22_port, S => q_2_2_22_port, Co => 
                           q_2_3_23_port);
   FA_C_1_3_23 : FA_533 port map( A => q_0_3_23_port, B => q_0_4_23_port, Ci =>
                           q_0_5_23_port, S => q_2_2_23_port, Co => 
                           q_2_3_24_port);
   FA_C_1_3_24 : FA_532 port map( A => q_0_4_24_port, B => q_0_5_24_port, Ci =>
                           q_0_6_24_port, S => n185, Co => q_2_3_25_port);
   FA_C_1_3_25 : FA_531 port map( A => q_0_3_25_port, B => q_0_4_25_port, Ci =>
                           q_0_5_25_port, S => q_2_2_25_port, Co => 
                           q_2_3_26_port);
   FA_C_1_3_26 : FA_530 port map( A => q_0_5_26_port, B => q_0_6_26_port, Ci =>
                           q_0_7_26_port, S => q_2_2_26_port, Co => 
                           q_2_3_27_port);
   FA_C_1_3_27 : FA_529 port map( A => q_1_3_27_port, B => q_0_5_27_port, Ci =>
                           q_0_6_27_port, S => q_2_2_27_port, Co => 
                           q_2_3_28_port);
   FA_C_1_3_28 : FA_528 port map( A => q_1_3_28_port, B => q_1_4_28_port, Ci =>
                           q_0_8_28_port, S => q_2_2_28_port, Co => 
                           q_2_3_29_port);
   FA_C_1_3_29 : FA_527 port map( A => q_1_3_29_port, B => q_1_4_29_port, Ci =>
                           q_1_5_29_port, S => q_2_2_29_port, Co => 
                           q_2_3_30_port);
   FA_C_1_3_30 : FA_526 port map( A => n190, B => q_1_4_30_port, Ci => 
                           q_1_5_30_port, S => q_2_2_30_port, Co => 
                           q_2_3_31_port);
   FA_C_1_3_31 : FA_525 port map( A => q_1_3_31_port, B => q_1_4_31_port, Ci =>
                           q_1_5_31_port, S => q_2_2_31_port, Co => 
                           q_2_3_32_port, clk => clk);
   FA_C_1_3_32 : FA_524 port map( A => q_1_3_32_port, B => q_1_4_32_port, Ci =>
                           q_1_5_32_port, S => q_2_2_32_port, Co => 
                           q_2_3_33_port);
   FA_C_1_3_33 : FA_523 port map( A => q_1_3_33_port, B => q_1_4_33_port, Ci =>
                           q_1_5_33_port, S => q_2_2_33_port, Co => 
                           q_2_3_34_port);
   FA_C_1_3_34 : FA_522 port map( A => q_1_3_34_port, B => q_1_4_34_port, Ci =>
                           q_1_5_34_port, S => q_2_2_34_port, Co => 
                           q_2_3_35_port);
   FA_C_1_3_35 : FA_521 port map( A => q_1_3_35_port, B => q_1_4_35_port, Ci =>
                           n184, S => q_2_2_35_port, Co => q_2_3_36_port);
   FA_C_1_3_36 : FA_520 port map( A => q_1_3_36_port, B => q_1_4_36_port, Ci =>
                           q_1_5_36_port, S => q_2_2_36_port, Co => 
                           q_2_3_37_port);
   FA_C_1_3_37 : FA_519 port map( A => q_1_3_37_port, B => q_1_4_37_port, Ci =>
                           q_1_5_37_port, S => q_2_2_37_port, Co => 
                           q_2_3_38_port, clk => clk);
   FA_C_1_3_38 : FA_518 port map( A => q_1_3_38_port, B => q_1_4_38_port, Ci =>
                           q_1_5_38_port, S => q_2_2_38_port, Co => 
                           q_2_3_39_port);
   FA_C_1_3_39 : FA_517 port map( A => q_1_3_39_port, B => q_1_4_39_port, Ci =>
                           q_0_6_39_port, S => q_2_2_39_port, Co => 
                           q_2_3_40_port);
   FA_C_1_3_40 : FA_516 port map( A => q_1_3_40_port, B => q_0_5_40_port, Ci =>
                           q_0_6_40_port, S => q_2_2_40_port, Co => 
                           q_2_3_41_port);
   FA_C_1_3_41 : FA_515 port map( A => q_0_3_41_port, B => q_0_4_41_port, Ci =>
                           q_0_5_41_port, S => q_2_2_41_port, Co => 
                           q_2_3_42_port);
   FA_C_1_3_42 : FA_514 port map( A => q_0_3_42_port, B => q_0_4_42_port, Ci =>
                           q_0_5_42_port, S => q_2_2_42_port, Co => 
                           q_2_3_43_port);
   FA_C_1_3_43 : FA_513 port map( A => q_0_2_43_port, B => q_0_3_43_port, Ci =>
                           q_0_4_43_port, S => q_2_2_43_port, Co => 
                           q_2_3_44_port);
   FA_C_1_3_44 : FA_512 port map( A => q_0_3_44_port, B => q_0_4_44_port, Ci =>
                           q_0_5_44_port, S => q_2_2_44_port, Co => 
                           q_2_3_45_port);
   FA_C_1_3_45 : FA_511 port map( A => q_0_3_45_port, B => q_0_4_45_port, Ci =>
                           q_0_5_45_port, S => q_2_2_45_port, Co => 
                           q_2_3_46_port);
   FA_C_1_3_46 : FA_510 port map( A => q_0_3_46_port, B => q_0_4_46_port, Ci =>
                           q_0_5_46_port, S => q_2_2_46_port, Co => 
                           q_2_3_47_port);
   FA_C_1_3_47 : FA_509 port map( A => q_0_3_47_port, B => q_0_4_47_port, Ci =>
                           q_0_5_47_port, S => q_2_2_47_port, Co => n_2383);
   HA_R_1_6_20 : HA_26 port map( A => q_0_6_20_port, B => q_0_7_20_port, S => 
                           n186, C => q_2_5_21_port);
   HA_R_1_6_21 : HA_25 port map( A => q_0_6_21_port, B => q_0_7_21_port, S => 
                           n188, C => q_2_5_22_port);
   FA_C_1_6_22 : FA_508 port map( A => q_0_6_22_port, B => q_0_7_22_port, Ci =>
                           q_0_8_22_port, S => q_2_4_22_port, Co => 
                           q_2_5_23_port);
   FA_C_1_6_23 : FA_507 port map( A => q_0_6_23_port, B => q_0_7_23_port, Ci =>
                           q_0_8_23_port, S => q_2_4_23_port, Co => 
                           q_2_5_24_port);
   FA_C_1_6_24 : FA_506 port map( A => q_0_7_24_port, B => q_0_8_24_port, Ci =>
                           q_0_9_24_port, S => q_2_4_24_port, Co => 
                           q_2_5_25_port);
   FA_C_1_6_25 : FA_505 port map( A => q_0_6_25_port, B => q_0_7_25_port, Ci =>
                           q_0_8_25_port, S => q_2_4_25_port, Co => 
                           q_2_5_26_port);
   FA_C_1_6_26 : FA_504 port map( A => q_0_8_26_port, B => q_0_9_26_port, Ci =>
                           q_0_10_26_port, S => q_2_4_26_port, Co => 
                           q_2_5_27_port);
   FA_C_1_6_27 : FA_503 port map( A => q_0_7_27_port, B => q_0_8_27_port, Ci =>
                           q_0_9_27_port, S => q_2_4_27_port, Co => 
                           q_2_5_28_port);
   FA_C_1_6_28 : FA_502 port map( A => q_0_9_28_port, B => q_0_10_28_port, Ci 
                           => q_0_11_28_port, S => q_2_4_28_port, Co => 
                           q_2_5_29_port);
   FA_C_1_6_29 : FA_501 port map( A => q_0_8_29_port, B => q_0_9_29_port, Ci =>
                           q_0_10_29_port, S => q_2_4_29_port, Co => 
                           q_2_5_30_port);
   FA_C_1_6_30 : FA_500 port map( A => n189, B => q_0_11_30_port, Ci => 
                           q_0_12_30_port, S => q_2_4_30_port, Co => 
                           q_2_5_31_port);
   FA_C_1_6_31 : FA_499 port map( A => q_1_6_31_port, B => q_1_7_31_port, Ci =>
                           q_0_11_31_port, S => q_2_4_31_port, Co => 
                           q_2_5_32_port);
   FA_C_1_6_32 : FA_498 port map( A => q_1_6_32_port, B => q_1_7_32_port, Ci =>
                           q_0_12_32_port, S => q_2_4_32_port, Co => 
                           q_2_5_33_port);
   FA_C_1_6_33 : FA_497 port map( A => q_1_6_33_port, B => q_1_7_33_port, Ci =>
                           q_0_12_33_port, S => q_2_4_33_port, Co => 
                           q_2_5_34_port, clk => clk);
   FA_C_1_6_34 : FA_496 port map( A => q_1_6_34_port, B => q_1_7_34_port, Ci =>
                           q_0_12_34_port, S => q_2_4_34_port, Co => 
                           q_2_5_35_port, clk => clk);
   FA_C_1_6_35 : FA_495 port map( A => q_1_6_35_port, B => q_1_7_35_port, Ci =>
                           q_0_12_35_port, S => q_2_4_35_port, Co => 
                           q_2_5_36_port);
   FA_C_1_6_36 : FA_494 port map( A => q_1_6_36_port, B => n179, Ci => 
                           q_0_11_36_port, S => q_2_4_36_port, Co => 
                           q_2_5_37_port);
   FA_C_1_6_37 : FA_493 port map( A => q_1_6_37_port, B => q_0_9_37_port, Ci =>
                           q_0_10_37_port, S => q_2_4_37_port, Co => 
                           q_2_5_38_port);
   FA_C_1_6_38 : FA_492 port map( A => q_0_8_38_port, B => q_0_9_38_port, Ci =>
                           q_0_10_38_port, S => q_2_4_38_port, Co => 
                           q_2_5_39_port);
   FA_C_1_6_39 : FA_491 port map( A => q_0_7_39_port, B => n191, Ci => 
                           q_0_9_39_port, S => q_2_4_39_port, Co => 
                           q_2_5_40_port);
   FA_C_1_6_40 : FA_490 port map( A => q_0_7_40_port, B => q_0_8_40_port, Ci =>
                           q_0_9_40_port, S => q_2_4_40_port, Co => 
                           q_2_5_41_port);
   FA_C_1_6_41 : FA_489 port map( A => q_0_6_41_port, B => q_0_7_41_port, Ci =>
                           q_0_8_41_port, S => q_2_4_41_port, Co => 
                           q_2_5_42_port);
   FA_C_1_6_42 : FA_488 port map( A => q_0_6_42_port, B => q_0_7_42_port, Ci =>
                           q_0_8_42_port, S => q_2_4_42_port, Co => 
                           q_2_5_43_port);
   FA_C_1_6_43 : FA_487 port map( A => q_0_5_43_port, B => q_0_6_43_port, Ci =>
                           q_0_7_43_port, S => q_2_4_43_port, Co => 
                           q_2_5_44_port);
   FA_C_1_6_44 : FA_486 port map( A => q_0_6_44_port, B => q_0_7_44_port, Ci =>
                           q_0_8_44_port, S => q_2_4_44_port, Co => 
                           q_2_5_45_port);
   FA_C_1_6_45 : FA_485 port map( A => q_0_6_45_port, B => q_0_7_45_port, Ci =>
                           q_0_8_45_port, S => q_2_4_45_port, Co => 
                           q_2_5_46_port);
   HA_L_1_6_46 : HA_24 port map( A => q_0_6_46_port, B => q_0_7_46_port, S => 
                           q_2_4_46_port, C => q_2_4_47_port);
   HA_R_1_9_22 : HA_23 port map( A => q_0_9_22_port, B => q_0_10_22_port, S => 
                           q_2_6_22_port, C => q_2_7_23_port);
   HA_R_1_9_23 : HA_22 port map( A => q_0_9_23_port, B => q_0_10_23_port, S => 
                           q_2_6_23_port, C => q_2_7_24_port);
   FA_C_1_9_24 : FA_484 port map( A => q_0_10_24_port, B => q_0_11_24_port, Ci 
                           => q_0_12_24_port, S => q_2_6_24_port, Co => 
                           q_2_7_25_port);
   FA_C_1_9_25 : FA_483 port map( A => q_0_9_25_port, B => q_0_10_25_port, Ci 
                           => q_0_11_25_port, S => q_2_6_25_port, Co => 
                           q_2_7_26_port);
   FA_C_1_9_26 : FA_482 port map( A => q_0_11_26_port, B => q_0_12_26_port, Ci 
                           => q_0_13_26_port, S => q_2_6_26_port, Co => 
                           q_2_7_27_port);
   FA_C_1_9_27 : FA_481 port map( A => q_0_10_27_port, B => q_0_11_27_port, Ci 
                           => q_0_12_27_port, S => q_2_6_27_port, Co => 
                           q_2_7_28_port);
   FA_C_1_9_28 : FA_480 port map( A => q_0_12_28_port, B => q_0_13_28_port, Ci 
                           => q_0_14_28_port, S => q_2_6_28_port, Co => 
                           q_2_7_29_port);
   FA_C_1_9_29 : FA_479 port map( A => q_0_11_29_port, B => q_0_12_29_port, Ci 
                           => q_0_13_29_port, S => n180, Co => q_2_7_30_port);
   FA_C_1_9_30 : FA_478 port map( A => q_0_13_30_port, B => q_0_14_30_port, Ci 
                           => net102771, S => q_2_6_30_port, clk => clk, Co_BAR
                           => q_2_7_31_port);
   FA_C_1_9_31 : FA_477 port map( A => q_0_12_31_port, B => q_0_13_31_port, Ci 
                           => q_0_14_31_port, S => q_2_6_31_port, Co => 
                           q_2_7_32_port);
   FA_C_1_9_32 : FA_476 port map( Ci => net102770, Co => q_2_7_33_port, B_BAR 
                           => q_0_14_32_port, A_BAR => q_0_13_32_port, S_BAR =>
                           q_2_6_32_port);
   FA_C_1_9_42 : FA_466 port map( B => net102768, Ci => net102769, Co => n_2384
                           , A_BAR => q_0_9_42_port, S_BAR => q_2_6_42_port);
   FA_C_1_9_43 : FA_465 port map( A => q_0_8_43_port, B => net102766, Ci => 
                           net102767, Co => n_2385, clk => clk, S_BAR => 
                           q_2_6_43_port);
   HA_L_1_9_44 : HA_21 port map( B => net102765, C => n_2386, S_BAR => 
                           q_2_6_44_port, A_BAR => q_0_9_44_port);
   HA_R_2_0_10 : HA_20 port map( A => q_0_0_10_port, B => q_0_1_10_port, S => 
                           n187, C => q_3_1_11_port);
   HA_R_2_0_11 : HA_19 port map( A => q_0_0_11_port, B => q_0_1_11_port, S => 
                           q_3_0_11_port, C => q_3_1_12_port);
   FA_C_2_0_12 : FA_464 port map( A => q_0_0_12_port, B => q_0_1_12_port, Ci =>
                           q_0_2_12_port, S => n183, Co => q_3_1_13_port);
   FA_C_2_0_13 : FA_463 port map( A => q_0_0_13_port, B => q_0_1_13_port, Ci =>
                           q_0_2_13_port, S => q_3_0_13_port, Co => 
                           q_3_1_14_port);
   FA_C_2_0_14 : FA_462 port map( A => q_0_0_14_port, B => q_0_1_14_port, Ci =>
                           q_0_2_14_port, S => q_3_0_14_port, Co => 
                           q_3_1_15_port);
   FA_C_2_0_15 : FA_461 port map( A => q_0_0_15_port, B => q_0_1_15_port, Ci =>
                           q_0_2_15_port, S => q_3_0_15_port, Co => 
                           q_3_1_16_port);
   FA_C_2_0_16 : FA_460 port map( A => q_2_0_16_port, B => q_0_2_16_port, Ci =>
                           q_0_3_16_port, S => q_3_0_16_port, Co => 
                           q_3_1_17_port);
   FA_C_2_0_17 : FA_459 port map( A => q_2_0_17_port, B => q_2_1_17_port, Ci =>
                           q_0_2_17_port, S => q_3_0_17_port, Co => 
                           q_3_1_18_port);
   FA_C_2_0_18 : FA_458 port map( A => q_2_0_18_port, B => q_2_1_18_port, Ci =>
                           q_2_2_18_port, S => q_3_0_18_port, Co => 
                           q_3_1_19_port);
   FA_C_2_0_19 : FA_457 port map( A => q_2_0_19_port, B => q_2_1_19_port, Ci =>
                           q_2_2_19_port, S => q_3_0_19_port, Co => 
                           q_3_1_20_port, clk => clk);
   FA_C_2_0_20 : FA_456 port map( A => q_2_0_20_port, B => q_2_1_20_port, Ci =>
                           q_2_2_20_port, S => q_3_0_20_port, Co => 
                           q_3_1_21_port, clk => clk);
   FA_C_2_0_21 : FA_455 port map( A => q_2_0_21_port, B => q_2_1_21_port, Ci =>
                           q_2_2_21_port, S => q_3_0_21_port, Co => 
                           q_3_1_22_port);
   FA_C_2_0_22 : FA_454 port map( A => q_2_0_22_port, B => q_2_1_22_port, Ci =>
                           q_2_2_22_port, S => q_3_0_22_port, Co => 
                           q_3_1_23_port);
   FA_C_2_0_23 : FA_453 port map( A => q_2_0_23_port, B => q_2_1_23_port, Ci =>
                           q_2_2_23_port, S => q_3_0_23_port, Co => 
                           q_3_1_24_port);
   FA_C_2_0_24 : FA_452 port map( A => q_2_0_24_port, B => q_2_1_24_port, Ci =>
                           n185, S => q_3_0_24_port, Co => q_3_1_25_port);
   FA_C_2_0_25 : FA_451 port map( A => q_2_0_25_port, B => q_2_1_25_port, Ci =>
                           q_2_2_25_port, S => q_3_0_25_port, Co => 
                           q_3_1_26_port, clk => clk);
   FA_C_2_0_26 : FA_450 port map( A => q_2_0_26_port, B => q_2_1_26_port, Ci =>
                           q_2_2_26_port, S => n201, Co => q_3_1_27_port, clk 
                           => clk);
   FA_C_2_0_27 : FA_449 port map( A => q_2_0_27_port, B => q_2_1_27_port, Ci =>
                           q_2_2_27_port, S => n196, Co => q_3_1_28_port, clk 
                           => clk);
   FA_C_2_0_28 : FA_448 port map( A => q_2_0_28_port, B => q_2_1_28_port, Ci =>
                           q_2_2_28_port, S => q_3_0_28_port, Co => 
                           q_3_1_29_port, clk => clk);
   FA_C_2_0_29 : FA_447 port map( A => q_2_0_29_port, B => q_2_1_29_port, Ci =>
                           q_2_2_29_port, S => q_3_0_29_port, Co => 
                           q_3_1_30_port, clk => clk);
   FA_C_2_0_30 : FA_446 port map( A => q_2_0_30_port, B => q_2_1_30_port, Ci =>
                           q_2_2_30_port, S => q_3_0_30_port, Co => 
                           q_3_1_31_port, clk => clk);
   FA_C_2_0_31 : FA_445 port map( A => q_2_0_31_port, B => q_2_1_31_port, Ci =>
                           q_2_2_31_port, S => q_3_0_31_port, Co => 
                           q_3_1_32_port, clk => clk);
   FA_C_2_0_32 : FA_444 port map( A => q_2_0_32_port, B => q_2_1_32_port, Ci =>
                           q_2_2_32_port, S => q_3_0_32_port, Co => 
                           q_3_1_33_port, clk => clk);
   FA_C_2_0_33 : FA_443 port map( A => q_2_0_33_port, B => q_2_1_33_port, Ci =>
                           q_2_2_33_port, S => q_3_0_33_port, Co => 
                           q_3_1_34_port, clk => clk);
   FA_C_2_0_34 : FA_442 port map( A => q_2_0_34_port, B => q_2_1_34_port, Ci =>
                           q_2_2_34_port, S => q_3_0_34_port, Co => 
                           q_3_1_35_port, clk => clk);
   FA_C_2_0_35 : FA_441 port map( A => q_2_0_35_port, B => q_2_1_35_port, Ci =>
                           q_2_2_35_port, S => q_3_0_35_port, Co => 
                           q_3_1_36_port, clk => clk);
   FA_C_2_0_36 : FA_440 port map( A => q_2_0_36_port, B => q_2_1_36_port, Ci =>
                           q_2_2_36_port, S => q_3_0_36_port, Co => 
                           q_3_1_37_port, clk => clk);
   FA_C_2_0_37 : FA_439 port map( A => q_2_0_37_port, B => q_2_1_37_port, Ci =>
                           q_2_2_37_port, S => q_3_0_37_port, Co => 
                           q_3_1_38_port, clk => clk);
   FA_C_2_0_38 : FA_438 port map( A => q_2_0_38_port, B => q_2_1_38_port, Ci =>
                           q_2_2_38_port, S => q_3_0_38_port, Co => 
                           q_3_1_39_port, clk => clk);
   FA_C_2_0_39 : FA_437 port map( A => q_2_0_39_port, B => q_2_1_39_port, Ci =>
                           q_2_2_39_port, S => q_3_0_39_port, Co => 
                           q_3_1_40_port, clk => clk);
   FA_C_2_0_40 : FA_436 port map( A => q_2_0_40_port, B => q_2_1_40_port, Ci =>
                           q_2_2_40_port, S => q_3_0_40_port, Co => 
                           q_3_1_41_port, clk => clk);
   FA_C_2_0_41 : FA_435 port map( A => q_2_0_41_port, B => q_2_1_41_port, Ci =>
                           q_2_2_41_port, S => q_3_0_41_port, Co => 
                           q_3_1_42_port, clk => clk);
   FA_C_2_0_42 : FA_434 port map( A => q_2_0_42_port, B => q_2_1_42_port, Ci =>
                           q_2_2_42_port, S => q_3_0_42_port, Co => 
                           q_3_1_43_port, clk => clk);
   FA_C_2_0_43 : FA_433 port map( A => q_2_0_43_port, B => q_2_1_43_port, Ci =>
                           q_2_2_43_port, S => q_3_0_43_port, Co => 
                           q_3_1_44_port, clk => clk);
   FA_C_2_0_44 : FA_432 port map( A => q_2_0_44_port, B => q_2_1_44_port, Ci =>
                           q_2_2_44_port, S => q_3_0_44_port, Co => 
                           q_3_1_45_port, clk => clk);
   FA_C_2_0_45 : FA_431 port map( A => q_2_0_45_port, B => q_2_1_45_port, Ci =>
                           q_2_2_45_port, S => q_3_0_45_port, Co => 
                           q_3_1_46_port);
   FA_C_2_0_46 : FA_430 port map( A => q_2_0_46_port, B => q_2_1_46_port, Ci =>
                           q_2_2_46_port, S => q_3_0_46_port, Co => 
                           q_3_1_47_port);
   FA_C_2_0_47 : FA_429 port map( A => q_2_0_47_port, B => q_2_1_47_port, Ci =>
                           q_2_2_47_port, S => q_3_0_47_port, Co => n_2387, clk
                           => clk);
   HA_R_2_3_12 : HA_17 port map( A => q_0_3_12_port, B => q_0_4_12_port, S => 
                           q_3_2_12_port, C => q_3_3_13_port);
   HA_R_2_3_13 : HA_16 port map( A => q_0_3_13_port, B => q_0_4_13_port, S => 
                           q_3_2_13_port, C => q_3_3_14_port);
   FA_C_2_3_14 : FA_420 port map( A => q_0_3_14_port, B => q_0_4_14_port, Ci =>
                           q_0_5_14_port, S => q_3_2_14_port, Co => 
                           q_3_3_15_port);
   FA_C_2_3_15 : FA_419 port map( A => q_0_3_15_port, B => q_0_4_15_port, Ci =>
                           q_0_5_15_port, S => q_3_2_15_port, Co => 
                           q_3_3_16_port);
   FA_C_2_3_16 : FA_418 port map( A => q_0_4_16_port, B => q_0_5_16_port, Ci =>
                           q_0_6_16_port, S => q_3_2_16_port, Co => 
                           q_3_3_17_port);
   FA_C_2_3_17 : FA_417 port map( A => q_0_3_17_port, B => q_0_4_17_port, Ci =>
                           q_0_5_17_port, S => q_3_2_17_port, Co => 
                           q_3_3_18_port);
   FA_C_2_3_18 : FA_416 port map( A => q_0_5_18_port, B => q_0_6_18_port, Ci =>
                           q_0_7_18_port, S => q_3_2_18_port, Co => 
                           q_3_3_19_port);
   FA_C_2_3_19 : FA_415 port map( A => q_2_3_19_port, B => q_0_5_19_port, Ci =>
                           q_0_6_19_port, S => q_3_2_19_port, Co => 
                           q_3_3_20_port);
   FA_C_2_3_20 : FA_414 port map( A => q_2_3_20_port, B => n186, Ci => 
                           q_0_8_20_port, S => q_3_2_20_port, Co => 
                           q_3_3_21_port);
   FA_C_2_3_21 : FA_413 port map( A => q_2_3_21_port, B => n188, Ci => 
                           q_2_5_21_port, S => q_3_2_21_port, Co => 
                           q_3_3_22_port);
   FA_C_2_3_22 : FA_412 port map( A => q_2_3_22_port, B => q_2_4_22_port, Ci =>
                           q_2_5_22_port, S => q_3_2_22_port, Co => 
                           q_3_3_23_port, clk => clk);
   FA_C_2_3_23 : FA_411 port map( A => q_2_3_23_port, B => q_2_4_23_port, Ci =>
                           q_2_5_23_port, S => q_3_2_23_port, Co => 
                           q_3_3_24_port);
   FA_C_2_3_24 : FA_410 port map( A => q_2_3_24_port, B => q_2_4_24_port, Ci =>
                           q_2_5_24_port, S => q_3_2_24_port, Co => 
                           q_3_3_25_port);
   FA_C_2_3_25 : FA_409 port map( A => q_2_3_25_port, B => q_2_4_25_port, Ci =>
                           q_2_5_25_port, S => q_3_2_25_port, Co => 
                           q_3_3_26_port);
   FA_C_2_3_26 : FA_408 port map( A => q_2_3_26_port, B => q_2_4_26_port, Ci =>
                           q_2_5_26_port, S => q_3_2_26_port, Co => 
                           q_3_3_27_port, clk => clk);
   FA_C_2_3_27 : FA_407 port map( A => q_2_3_27_port, B => q_2_4_27_port, Ci =>
                           q_2_5_27_port, S => q_3_2_27_port, Co => 
                           q_3_3_28_port, clk => clk);
   FA_C_2_3_28 : FA_406 port map( A => q_2_3_28_port, B => q_2_4_28_port, Ci =>
                           q_2_5_28_port, S => q_3_2_28_port, Co => 
                           q_3_3_29_port, clk => clk);
   FA_C_2_3_29 : FA_405 port map( A => q_2_3_29_port, B => q_2_4_29_port, Ci =>
                           q_2_5_29_port, S => q_3_2_29_port, Co => 
                           q_3_3_30_port, clk => clk);
   FA_C_2_3_30 : FA_404 port map( A => q_2_3_30_port, B => q_2_4_30_port, Ci =>
                           q_2_5_30_port, S => q_3_2_30_port, Co => 
                           q_3_3_31_port, clk => clk);
   FA_C_2_3_31 : FA_403 port map( A => q_2_3_31_port, B => q_2_4_31_port, Ci =>
                           q_2_5_31_port, S => q_3_2_31_port, Co => 
                           q_3_3_32_port, clk => clk);
   FA_C_2_3_32 : FA_402 port map( A => q_2_3_32_port, B => q_2_4_32_port, Ci =>
                           q_2_5_32_port, S => q_3_2_32_port, Co => 
                           q_3_3_33_port, clk => clk);
   FA_C_2_3_33 : FA_401 port map( A => q_2_3_33_port, B => q_2_4_33_port, Ci =>
                           q_2_5_33_port, S => q_3_2_33_port, Co => 
                           q_3_3_34_port, clk => clk);
   FA_C_2_3_34 : FA_400 port map( A => q_2_3_34_port, B => q_2_4_34_port, Ci =>
                           q_2_5_34_port, S => q_3_2_34_port, Co => 
                           q_3_3_35_port, clk => clk);
   FA_C_2_3_35 : FA_399 port map( A => q_2_3_35_port, B => q_2_4_35_port, Ci =>
                           q_2_5_35_port, S => q_3_2_35_port, Co => 
                           q_3_3_36_port, clk => clk);
   FA_C_2_3_36 : FA_398 port map( A => q_2_3_36_port, B => q_2_4_36_port, Ci =>
                           q_2_5_36_port, S => q_3_2_36_port, Co => 
                           q_3_3_37_port, clk => clk);
   FA_C_2_3_37 : FA_397 port map( A => q_2_3_37_port, B => q_2_4_37_port, Ci =>
                           q_2_5_37_port, S => q_3_2_37_port, Co => 
                           q_3_3_38_port, clk => clk);
   FA_C_2_3_38 : FA_396 port map( A => q_2_3_38_port, B => q_2_4_38_port, Ci =>
                           q_2_5_38_port, S => q_3_2_38_port, Co => 
                           q_3_3_39_port, clk => clk);
   FA_C_2_3_39 : FA_395 port map( A => q_2_3_39_port, B => q_2_4_39_port, Ci =>
                           q_2_5_39_port, S => q_3_2_39_port, Co => 
                           q_3_3_40_port, clk => clk);
   FA_C_2_3_40 : FA_394 port map( A => q_2_3_40_port, B => q_2_4_40_port, Ci =>
                           q_2_5_40_port, S => q_3_2_40_port, Co => 
                           q_3_3_41_port, clk => clk);
   FA_C_2_3_41 : FA_393 port map( A => q_2_3_41_port, B => q_2_4_41_port, Ci =>
                           q_2_5_41_port, S => q_3_2_41_port, Co => 
                           q_3_3_42_port, clk => clk);
   FA_C_2_3_42 : FA_392 port map( A => q_2_3_42_port, B => q_2_4_42_port, Ci =>
                           q_2_5_42_port, S => q_3_2_42_port, Co => 
                           q_3_3_43_port, clk => clk);
   FA_C_2_3_43 : FA_391 port map( A => q_2_3_43_port, B => q_2_4_43_port, Ci =>
                           q_2_5_43_port, S => q_3_2_43_port, Co => 
                           q_3_3_44_port, clk => clk);
   FA_C_2_3_44 : FA_390 port map( A => q_2_3_44_port, B => q_2_4_44_port, Ci =>
                           q_2_5_44_port, S => q_3_2_44_port, Co => 
                           q_3_3_45_port, clk => clk);
   FA_C_2_3_45 : FA_389 port map( A => q_2_3_45_port, B => q_2_4_45_port, Ci =>
                           q_2_5_45_port, S => q_3_2_45_port, Co => 
                           q_3_3_46_port, clk => clk);
   FA_C_2_3_46 : FA_388 port map( A => q_2_3_46_port, B => q_2_4_46_port, Ci =>
                           q_2_5_46_port, S => q_3_2_46_port, Co => 
                           q_3_3_47_port, clk => clk);
   FA_C_2_3_47 : FA_387 port map( A => q_2_3_47_port, B => q_2_4_47_port, Ci =>
                           q_0_6_47_port, S => q_3_2_47_port, Co => n_2388);
   HA_R_2_6_14 : HA_14 port map( A => q_0_6_14_port, B => q_0_7_14_port, S => 
                           n192, C => q_3_5_15_port);
   HA_R_2_6_15 : HA_13 port map( A => q_0_6_15_port, B => q_0_7_15_port, S => 
                           q_3_4_15_port, C => q_3_5_16_port);
   FA_C_2_6_16 : FA_380 port map( A => q_0_7_16_port, B => q_0_8_16_port, Ci =>
                           B(17), S => q_3_4_16_port, Co => q_3_5_17_port);
   FA_C_2_6_17 : FA_379 port map( A => q_0_6_17_port, B => q_0_7_17_port, Ci =>
                           q_0_8_17_port, S => q_3_4_17_port, Co => 
                           q_3_5_18_port);
   FA_C_2_6_18 : FA_378 port map( A => q_0_8_18_port, B => q_0_9_18_port, Ci =>
                           B(19), S => q_3_4_18_port, Co => q_3_5_19_port);
   FA_C_2_6_19 : FA_377 port map( A => q_0_7_19_port, B => q_0_8_19_port, Ci =>
                           q_0_9_19_port, S => q_3_4_19_port, Co => 
                           q_3_5_20_port);
   FA_C_2_6_20 : FA_376 port map( A => q_0_9_20_port, B => q_0_10_20_port, Ci 
                           => B(21), S => q_3_4_20_port, Co => q_3_5_21_port);
   FA_C_2_6_21 : FA_375 port map( A => q_0_8_21_port, B => q_0_9_21_port, Ci =>
                           q_0_10_21_port, S => q_3_4_21_port, Co => 
                           q_3_5_22_port);
   FA_C_2_6_22 : FA_374 port map( A => q_2_6_22_port, B => q_0_11_22_port, Ci 
                           => n2, S => q_3_4_22_port, Co => q_3_5_23_port);
   FA_C_2_6_23 : FA_373 port map( A => q_2_6_23_port, B => q_2_7_23_port, Ci =>
                           q_0_11_23_port, S => q_3_4_23_port, Co => 
                           q_3_5_24_port);
   FA_C_2_6_24 : FA_372 port map( A => q_2_6_24_port, B => q_2_7_24_port, Ci =>
                           n213, S => q_3_4_24_port, Co => q_3_5_25_port);
   FA_C_2_6_25 : FA_371 port map( A => q_2_6_25_port, B => q_2_7_25_port, Ci =>
                           q_0_12_25_port, S => q_3_4_25_port, Co => 
                           q_3_5_26_port, clk => clk);
   FA_C_2_6_26 : FA_370 port map( A => q_2_6_26_port, B => q_2_7_26_port, Ci =>
                           n211, S => q_3_4_26_port, Co => q_3_5_27_port, clk 
                           => clk);
   FA_C_2_6_27 : FA_369 port map( A => q_2_6_27_port, B => q_2_7_27_port, Ci =>
                           q_0_13_27_port, S => q_3_4_27_port, Co => 
                           q_3_5_28_port, clk => clk);
   FA_C_2_6_28 : FA_368 port map( A => q_2_6_28_port, B => q_2_7_28_port, Ci =>
                           n209, S => q_3_4_28_port, Co => q_3_5_29_port, clk 
                           => clk);
   FA_C_2_6_29 : FA_367 port map( A => n180, B => q_2_7_29_port, Ci => 
                           q_0_14_29_port, S => q_3_4_29_port, Co => 
                           q_3_5_30_port);
   FA_C_2_6_30 : FA_366 port map( A => q_2_6_30_port, B => q_2_7_30_port, Ci =>
                           n207, S => q_3_4_30_port, Co => q_3_5_31_port, clk 
                           => clk);
   FA_C_2_6_31 : FA_365 port map( A => q_2_6_31_port, Ci => net102764, S => 
                           q_3_4_31_port, Co => q_3_5_32_port, clk => clk, 
                           B_BAR => q_2_7_31_port);
   FA_C_2_6_32 : FA_364 port map( B => q_2_7_32_port, Ci => net102763, S => 
                           q_3_4_32_port, Co => q_3_5_33_port, clk => clk, 
                           A_BAR => q_2_6_32_port);
   FA_C_2_6_33 : FA_363 port map( A => net102761, B => q_2_7_33_port, Ci => 
                           net102762, S => q_3_4_33_port, Co => n_2389);
   FA_C_2_6_42 : FA_354 port map( B => net102759, Ci => net102760, Co => n_2390
                           , A_BAR => q_2_6_42_port, S_BAR => q_3_4_42_port);
   FA_C_2_6_43 : FA_353 port map( B => net102757, Ci => net102758, Co => n_2391
                           , A_BAR => q_2_6_43_port, S_BAR => q_3_4_43_port);
   FA_C_2_6_44 : FA_352 port map( B => net102755, Ci => net102756, Co => n_2392
                           , A_BAR => q_2_6_44_port, S_BAR => q_3_4_44_port);
   FA_C_2_6_46 : FA_350 port map( A => q_0_8_46_port, S => q_3_4_46_port, Co =>
                           q_3_5_47_port, clk => clk, Ci_BAR => q_0_10_46_port,
                           B_BAR => q_0_9_46_port);
   FA_C_2_6_47 : FA_349 port map( A => q_0_7_47_port, B => q_0_8_47_port, Ci =>
                           q_0_9_47_port, S => q_3_4_47_port, Co => n_2393);
   HA_R_3_0_6 : HA_11 port map( A => q_0_0_6_port, B => q_0_1_6_port, S => 
                           q_4_0_6_port, C => q_4_1_7_port);
   HA_R_3_0_7 : HA_10 port map( A => q_0_0_7_port, B => q_0_1_7_port, S => 
                           q_4_0_7_port, C => q_4_1_8_port);
   FA_C_3_0_8 : FA_344 port map( A => q_0_0_8_port, B => q_0_1_8_port, Ci => 
                           q_0_2_8_port, S => q_4_0_8_port, Co => q_4_1_9_port)
                           ;
   FA_C_3_0_9 : FA_343 port map( A => q_0_0_9_port, B => q_0_1_9_port, Ci => 
                           q_0_2_9_port, S => q_4_0_9_port, Co => q_4_1_10_port
                           );
   FA_C_3_0_10 : FA_342 port map( A => n187, B => q_0_2_10_port, Ci => 
                           q_0_3_10_port, S => q_4_0_10_port, Co => 
                           q_4_1_11_port);
   FA_C_3_0_11 : FA_341 port map( A => q_3_0_11_port, B => q_3_1_11_port, Ci =>
                           q_0_2_11_port, S => q_4_0_11_port, Co => 
                           q_4_1_12_port);
   FA_C_3_0_12 : FA_340 port map( A => n183, B => q_3_1_12_port, Ci => 
                           q_3_2_12_port, S => q_4_0_12_port, Co => 
                           q_4_1_13_port);
   FA_C_3_0_13 : FA_339 port map( A => q_3_0_13_port, B => q_3_1_13_port, Ci =>
                           q_3_2_13_port, S => q_4_0_13_port, Co => 
                           q_4_1_14_port, clk => clk);
   FA_C_3_0_14 : FA_338 port map( A => q_3_0_14_port, B => q_3_1_14_port, Ci =>
                           q_3_2_14_port, S => q_4_0_14_port, Co => 
                           q_4_1_15_port);
   FA_C_3_0_15 : FA_337 port map( A => q_3_0_15_port, B => q_3_1_15_port, Ci =>
                           q_3_2_15_port, S => q_4_0_15_port, Co => 
                           q_4_1_16_port);
   FA_C_3_0_16 : FA_336 port map( A => q_3_0_16_port, B => q_3_1_16_port, Ci =>
                           q_3_2_16_port, S => q_4_0_16_port, Co => 
                           q_4_1_17_port, clk => clk);
   FA_C_3_0_17 : FA_335 port map( A => q_3_0_17_port, B => q_3_1_17_port, Ci =>
                           q_3_2_17_port, S => q_4_0_17_port, Co => 
                           q_4_1_18_port, clk => clk);
   FA_C_3_0_18 : FA_334 port map( A => q_3_0_18_port, B => q_3_1_18_port, Ci =>
                           q_3_2_18_port, S => q_4_0_18_port, Co => 
                           q_4_1_19_port, clk => clk);
   FA_C_3_0_19 : FA_333 port map( A => q_3_0_19_port, B => q_3_1_19_port, Ci =>
                           q_3_2_19_port, S => q_4_0_19_port, Co => 
                           q_4_1_20_port, clk => clk);
   FA_C_3_0_20 : FA_332 port map( A => q_3_0_20_port, B => q_3_1_20_port, Ci =>
                           q_3_2_20_port, S => q_4_0_20_port, Co => 
                           q_4_1_21_port, clk => clk);
   FA_C_3_0_21 : FA_331 port map( A => q_3_0_21_port, B => q_3_1_21_port, Ci =>
                           q_3_2_21_port, S => q_4_0_21_port, Co => 
                           q_4_1_22_port, clk => clk);
   FA_C_3_0_22 : FA_330 port map( A => q_3_0_22_port, B => q_3_1_22_port, Ci =>
                           q_3_2_22_port, S => n199, Co => q_4_1_23_port, clk 
                           => clk);
   FA_C_3_0_23 : FA_329 port map( A => q_3_0_23_port, B => q_3_1_23_port, Ci =>
                           q_3_2_23_port, S => n195, Co => q_4_1_24_port, clk 
                           => clk);
   FA_C_3_0_24 : FA_328 port map( A => q_3_0_24_port, B => q_3_1_24_port, Ci =>
                           q_3_2_24_port, S => q_4_0_24_port, Co => 
                           q_4_1_25_port, clk => clk);
   FA_C_3_0_25 : FA_327 port map( A => q_3_0_25_port, B => q_3_1_25_port, Ci =>
                           q_3_2_25_port, S => n194, Co => q_4_1_26_port, clk 
                           => clk);
   FA_C_3_0_26 : FA_326 port map( A => n201, B => q_3_1_26_port, Ci => 
                           q_3_2_26_port, S => q_4_0_26_port, Co => 
                           q_4_1_27_port);
   FA_C_3_0_27 : FA_325 port map( A => n196, B => q_3_1_27_port, Ci => 
                           q_3_2_27_port, S => q_4_0_27_port, Co => 
                           q_4_1_28_port);
   FA_C_3_0_28 : FA_324 port map( A => q_3_0_28_port, B => q_3_1_28_port, Ci =>
                           q_3_2_28_port, S => q_4_0_28_port, Co => 
                           q_4_1_29_port);
   FA_C_3_0_29 : FA_323 port map( A => q_3_0_29_port, B => q_3_1_29_port, Ci =>
                           q_3_2_29_port, S => q_4_0_29_port, Co => 
                           q_4_1_30_port);
   FA_C_3_0_30 : FA_322 port map( A => q_3_0_30_port, B => q_3_1_30_port, Ci =>
                           q_3_2_30_port, S => q_4_0_30_port, Co => 
                           q_4_1_31_port);
   FA_C_3_0_31 : FA_321 port map( A => q_3_0_31_port, B => q_3_1_31_port, Ci =>
                           q_3_2_31_port, S => q_4_0_31_port, Co => 
                           q_4_1_32_port);
   FA_C_3_0_32 : FA_320 port map( A => q_3_0_32_port, B => q_3_1_32_port, Ci =>
                           q_3_2_32_port, S => q_4_0_32_port, Co => 
                           q_4_1_33_port);
   FA_C_3_0_33 : FA_319 port map( A => q_3_0_33_port, B => q_3_1_33_port, Ci =>
                           q_3_2_33_port, S => q_4_0_33_port, Co => 
                           q_4_1_34_port);
   FA_C_3_0_34 : FA_318 port map( A => q_3_0_34_port, B => q_3_1_34_port, Ci =>
                           q_3_2_34_port, S => q_4_0_34_port, Co => 
                           q_4_1_35_port);
   FA_C_3_0_35 : FA_317 port map( A => q_3_0_35_port, B => q_3_1_35_port, Ci =>
                           q_3_2_35_port, S => q_4_0_35_port, Co => 
                           q_4_1_36_port);
   FA_C_3_0_36 : FA_316 port map( A => q_3_0_36_port, B => q_3_1_36_port, Ci =>
                           q_3_2_36_port, S => q_4_0_36_port, Co => 
                           q_4_1_37_port);
   FA_C_3_0_37 : FA_315 port map( A => q_3_0_37_port, B => q_3_1_37_port, Ci =>
                           q_3_2_37_port, S => q_4_0_37_port, Co => 
                           q_4_1_38_port);
   FA_C_3_0_38 : FA_314 port map( A => q_3_0_38_port, B => q_3_1_38_port, Ci =>
                           q_3_2_38_port, S => q_4_0_38_port, Co => 
                           q_4_1_39_port);
   FA_C_3_0_39 : FA_313 port map( A => q_3_0_39_port, B => q_3_1_39_port, Ci =>
                           q_3_2_39_port, S => q_4_0_39_port, Co => 
                           q_4_1_40_port);
   FA_C_3_0_40 : FA_312 port map( A => q_3_0_40_port, B => q_3_1_40_port, Ci =>
                           q_3_2_40_port, S => q_4_0_40_port, Co => 
                           q_4_1_41_port);
   FA_C_3_0_41 : FA_311 port map( A => q_3_0_41_port, B => q_3_1_41_port, Ci =>
                           q_3_2_41_port, S => q_4_0_41_port, Co => 
                           q_4_1_42_port);
   FA_C_3_0_42 : FA_310 port map( A => q_3_0_42_port, B => q_3_1_42_port, Ci =>
                           q_3_2_42_port, S => q_4_0_42_port, Co => 
                           q_4_1_43_port);
   FA_C_3_0_43 : FA_309 port map( A => q_3_0_43_port, B => q_3_1_43_port, Ci =>
                           q_3_2_43_port, S => q_4_0_43_port, Co => 
                           q_4_1_44_port);
   FA_C_3_0_44 : FA_308 port map( A => q_3_0_44_port, B => q_3_1_44_port, Ci =>
                           q_3_2_44_port, S => q_4_0_44_port, Co => 
                           q_4_1_45_port, clk => clk);
   FA_C_3_0_45 : FA_307 port map( A => q_3_0_45_port, B => q_3_1_45_port, Ci =>
                           q_3_2_45_port, S => q_4_0_45_port, Co => 
                           q_4_1_46_port, clk => clk);
   FA_C_3_0_46 : FA_306 port map( A => q_3_0_46_port, B => q_3_1_46_port, Ci =>
                           q_3_2_46_port, S => q_4_0_46_port, Co => 
                           q_4_1_47_port, clk => clk);
   FA_C_3_0_47 : FA_305 port map( A => q_3_0_47_port, B => q_3_1_47_port, Ci =>
                           q_3_2_47_port, S => q_4_0_47_port, Co => n_2394, clk
                           => clk);
   HA_R_3_3_8 : HA_8 port map( A => q_0_3_8_port, B => q_0_4_8_port, S => 
                           q_4_2_8_port, C => q_5_2_9_port);
   HA_R_3_3_9 : HA_7 port map( A => q_0_3_9_port, B => q_0_4_9_port, S => 
                           q_4_2_9_port, C => q_5_2_10_port);
   FA_C_3_3_10 : FA_292 port map( A => q_0_4_10_port, B => q_0_5_10_port, Ci =>
                           B(11), S => q_4_2_10_port, Co => q_5_2_11_port);
   FA_C_3_3_11 : FA_291 port map( A => q_0_3_11_port, B => q_0_4_11_port, Ci =>
                           q_0_5_11_port, S => q_4_2_11_port, Co => 
                           q_5_2_12_port);
   FA_C_3_3_12 : FA_290 port map( A => q_0_5_12_port, B => q_0_6_12_port, S => 
                           q_4_2_12_port, Co => q_5_2_13_port, Ci => B(13));
   FA_C_3_3_13 : FA_289 port map( A => q_3_3_13_port, B => q_0_5_13_port, Ci =>
                           q_0_6_13_port, S => q_4_2_13_port, Co => 
                           q_5_2_14_port);
   FA_C_3_3_14 : FA_288 port map( A => q_3_3_14_port, B => n192, Ci => B(15), S
                           => q_4_2_14_port, Co => q_5_2_15_port);
   FA_C_3_3_15 : FA_287 port map( A => q_3_3_15_port, B => q_3_4_15_port, Ci =>
                           q_3_5_15_port, S => q_4_2_15_port, Co => 
                           q_5_2_16_port, clk => clk);
   FA_C_3_3_16 : FA_286 port map( A => q_3_3_16_port, B => q_3_4_16_port, Ci =>
                           q_3_5_16_port, S => q_4_2_16_port, Co => 
                           q_5_2_17_port, clk => clk);
   FA_C_3_3_17 : FA_285 port map( A => q_3_3_17_port, B => q_3_4_17_port, Ci =>
                           q_3_5_17_port, S => q_4_2_17_port, Co => 
                           q_5_2_18_port, clk => clk);
   FA_C_3_3_18 : FA_284 port map( A => q_3_3_18_port, B => q_3_4_18_port, Ci =>
                           q_3_5_18_port, S => q_4_2_18_port, Co => 
                           q_5_2_19_port, clk => clk);
   FA_C_3_3_19 : FA_283 port map( A => q_3_3_19_port, B => q_3_4_19_port, Ci =>
                           q_3_5_19_port, S => q_4_2_19_port, Co => 
                           q_5_2_20_port, clk => clk);
   FA_C_3_3_20 : FA_282 port map( A => q_3_3_20_port, B => q_3_4_20_port, Ci =>
                           q_3_5_20_port, S => n198, Co => q_5_2_21_port, clk 
                           => clk);
   FA_C_3_3_21 : FA_281 port map( A => q_3_3_21_port, B => q_3_4_21_port, Ci =>
                           q_3_5_21_port, S => q_4_2_21_port, Co => 
                           q_5_2_22_port, clk => clk);
   FA_C_3_3_22 : FA_280 port map( A => q_3_3_22_port, B => q_3_4_22_port, Ci =>
                           q_3_5_22_port, S => n197, Co => q_5_2_23_port, clk 
                           => clk);
   FA_C_3_3_23 : FA_279 port map( A => q_3_3_23_port, B => q_3_4_23_port, Ci =>
                           q_3_5_23_port, S => n200, Co => q_5_2_24_port, clk 
                           => clk);
   FA_C_3_3_24 : FA_278 port map( A => q_3_3_24_port, B => q_3_4_24_port, Ci =>
                           q_3_5_24_port, S => q_4_2_24_port, Co => 
                           q_5_2_25_port, clk => clk);
   FA_C_3_3_25 : FA_277 port map( A => q_3_3_25_port, B => q_3_4_25_port, Ci =>
                           q_3_5_25_port, S => q_4_2_25_port, Co => 
                           q_5_2_26_port, clk => clk);
   FA_C_3_3_26 : FA_276 port map( A => q_3_3_26_port, B => q_3_4_26_port, Ci =>
                           q_3_5_26_port, S => q_4_2_26_port, Co => 
                           q_5_2_27_port, clk => clk);
   FA_C_3_3_27 : FA_275 port map( A => q_3_3_27_port, B => q_3_4_27_port, Ci =>
                           q_3_5_27_port, S => q_4_2_27_port, Co => 
                           q_5_2_28_port, clk => clk);
   FA_C_3_3_28 : FA_274 port map( A => q_3_3_28_port, B => q_3_4_28_port, Ci =>
                           q_3_5_28_port, S => q_4_2_28_port, Co => 
                           q_5_2_29_port, clk => clk);
   FA_C_3_3_29 : FA_273 port map( A => q_3_3_29_port, B => q_3_4_29_port, Ci =>
                           q_3_5_29_port, S => q_4_2_29_port, Co => 
                           q_5_2_30_port, clk => clk);
   FA_C_3_3_30 : FA_272 port map( A => q_3_3_30_port, B => q_3_4_30_port, Ci =>
                           q_3_5_30_port, S => q_4_2_30_port, Co => 
                           q_5_2_31_port, clk => clk);
   FA_C_3_3_31 : FA_271 port map( A => q_3_3_31_port, B => q_3_4_31_port, Ci =>
                           q_3_5_31_port, S => q_4_2_31_port, Co => 
                           q_5_2_32_port);
   FA_C_3_3_32 : FA_270 port map( A => q_3_3_32_port, B => q_3_4_32_port, Ci =>
                           q_3_5_32_port, S => q_4_2_32_port, Co => 
                           q_5_2_33_port);
   FA_C_3_3_33 : FA_269 port map( A => q_3_3_33_port, B => q_3_4_33_port, Ci =>
                           q_3_5_33_port, S => q_4_2_33_port, Co => 
                           q_5_2_34_port);
   FA_C_3_3_34 : FA_268 port map( A => q_3_3_34_port, B => net102753, Ci => 
                           net102754, Co => n_2395, S => q_4_2_34_port);
   FA_C_3_3_35 : FA_267 port map( A => q_3_3_35_port, B => net102751, Ci => 
                           net102752, S => q_4_2_35_port, Co => n_2396);
   FA_C_3_3_36 : FA_266 port map( A => q_3_3_36_port, B => net102749, Ci => 
                           net102750, S => q_4_2_36_port, Co => n_2397);
   FA_C_3_3_37 : FA_265 port map( A => q_3_3_37_port, B => net102747, Ci => 
                           net102748, Co => n_2398, S => q_4_2_37_port);
   FA_C_3_3_38 : FA_264 port map( A => q_3_3_38_port, B => net102745, Ci => 
                           net102746, Co => n_2399, S => q_4_2_38_port);
   FA_C_3_3_39 : FA_263 port map( A => q_3_3_39_port, B => net102743, Ci => 
                           net102744, S => q_4_2_39_port, Co => n_2400);
   FA_C_3_3_40 : FA_262 port map( A => q_3_3_40_port, B => net102741, Ci => 
                           net102742, S => q_4_2_40_port, Co => n_2401);
   FA_C_3_3_41 : FA_261 port map( A => q_3_3_41_port, B => net102739, Ci => 
                           net102740, S => q_4_2_41_port, Co => n_2402);
   FA_C_3_3_42 : FA_260 port map( A => q_3_3_42_port, Ci => net102738, S => 
                           q_4_2_42_port, Co => q_5_2_43_port, B_BAR => 
                           q_3_4_42_port);
   FA_C_3_3_43 : FA_259 port map( A => q_3_3_43_port, Ci => net102737, S => 
                           q_4_2_43_port, Co => q_5_2_44_port, B_BAR => 
                           q_3_4_43_port);
   FA_C_3_3_44 : FA_258 port map( A => q_3_3_44_port, Ci => net102736, Co => 
                           q_5_2_45_port, B_BAR => q_3_4_44_port, S_BAR => 
                           q_4_2_44_port);
   FA_C_3_3_45 : FA_257 port map( A => q_3_3_45_port, B => net102734, Ci => 
                           net102735, Co => n_2403, S => q_4_2_45_port);
   FA_C_3_3_46 : FA_256 port map( A => q_3_3_46_port, B => q_3_4_46_port, Ci =>
                           net102733, Co => q_5_2_47_port, S_BAR => 
                           q_4_2_46_port);
   FA_C_3_3_47 : FA_255 port map( A => q_3_3_47_port, B => q_3_4_47_port, Ci =>
                           q_3_5_47_port, S => q_4_2_47_port, Co => n_2404, clk
                           => clk);
   HA_R_4_0_4 : HA_5 port map( A => q_0_0_4_port, B => q_0_1_4_port, S => 
                           q_5_0_4_port, C => q_5_1_5_port);
   HA_R_4_0_5 : HA_4 port map( A => q_0_0_5_port, B => q_0_1_5_port, S => 
                           q_5_0_5_port, C => q_5_1_6_port);
   FA_C_4_0_6 : FA_244 port map( A => q_4_0_6_port, B => q_0_2_6_port, Ci => 
                           q_0_3_6_port, S => q_5_0_6_port, Co => q_5_1_7_port)
                           ;
   FA_C_4_0_7 : FA_243 port map( A => q_4_0_7_port, B => q_4_1_7_port, Ci => 
                           q_0_2_7_port, S => q_5_0_7_port, Co => q_5_1_8_port)
                           ;
   FA_C_4_0_8 : FA_242 port map( A => q_4_0_8_port, B => q_4_1_8_port, Ci => 
                           q_4_2_8_port, S => q_5_0_8_port, Co => q_5_1_9_port,
                           clk => clk);
   FA_C_4_0_9 : FA_241 port map( A => q_4_0_9_port, B => q_4_1_9_port, Ci => 
                           q_4_2_9_port, S => q_5_0_9_port, Co => q_5_1_10_port
                           , clk => clk);
   FA_C_4_0_10 : FA_240 port map( A => q_4_0_10_port, B => q_4_1_10_port, Ci =>
                           q_4_2_10_port, S => q_5_0_10_port, Co => 
                           q_5_1_11_port, clk => clk);
   FA_C_4_0_11 : FA_239 port map( A => q_4_0_11_port, B => q_4_1_11_port, Ci =>
                           q_4_2_11_port, S => q_5_0_11_port, Co => 
                           q_5_1_12_port, clk => clk);
   FA_C_4_0_12 : FA_238 port map( A => q_4_0_12_port, B => q_4_1_12_port, Ci =>
                           q_4_2_12_port, S => q_5_0_12_port, Co => 
                           q_5_1_13_port, clk => clk);
   FA_C_4_0_13 : FA_237 port map( A => q_4_0_13_port, B => q_4_1_13_port, Ci =>
                           q_4_2_13_port, S => q_5_0_13_port, Co => 
                           q_5_1_14_port, clk => clk);
   FA_C_4_0_14 : FA_236 port map( A => q_4_0_14_port, B => q_4_1_14_port, Ci =>
                           q_4_2_14_port, S => q_5_0_14_port, Co => 
                           q_5_1_15_port, clk => clk);
   FA_C_4_0_15 : FA_235 port map( A => q_4_0_15_port, B => q_4_1_15_port, Ci =>
                           q_4_2_15_port, S => q_5_0_15_port, Co => 
                           q_5_1_16_port, clk => clk);
   FA_C_4_0_16 : FA_234 port map( A => q_4_0_16_port, B => q_4_1_16_port, Ci =>
                           q_4_2_16_port, S => n193, Co => q_5_1_17_port, clk 
                           => clk);
   FA_C_4_0_17 : FA_233 port map( A => q_4_0_17_port, B => q_4_1_17_port, Ci =>
                           q_4_2_17_port, S => q_5_0_17_port, Co => 
                           q_5_1_18_port, clk => clk);
   FA_C_4_0_18 : FA_232 port map( A => q_4_0_18_port, B => q_4_1_18_port, Ci =>
                           q_4_2_18_port, S => q_5_0_18_port, Co => 
                           q_5_1_19_port);
   FA_C_4_0_19 : FA_231 port map( A => q_4_0_19_port, B => q_4_1_19_port, Ci =>
                           q_4_2_19_port, S => q_5_0_19_port, Co => 
                           q_5_1_20_port);
   FA_C_4_0_20 : FA_230 port map( A => q_4_0_20_port, B => q_4_1_20_port, Ci =>
                           n198, S => q_5_0_20_port, Co => q_5_1_21_port);
   FA_C_4_0_21 : FA_229 port map( A => q_4_0_21_port, B => q_4_1_21_port, Ci =>
                           q_4_2_21_port, S => q_5_0_21_port, Co => 
                           q_5_1_22_port);
   FA_C_4_0_22 : FA_228 port map( A => n199, B => q_4_1_22_port, Ci => n197, S 
                           => q_5_0_22_port, Co => q_5_1_23_port);
   FA_C_4_0_23 : FA_227 port map( A => n195, B => q_4_1_23_port, Ci => n200, S 
                           => q_5_0_23_port, Co => q_5_1_24_port);
   FA_C_4_0_24 : FA_226 port map( A => q_4_0_24_port, B => q_4_1_24_port, Ci =>
                           q_4_2_24_port, S => q_5_0_24_port, Co => 
                           q_5_1_25_port);
   FA_C_4_0_25 : FA_225 port map( A => n194, B => q_4_1_25_port, Ci => 
                           q_4_2_25_port, S => q_5_0_25_port, Co => 
                           q_5_1_26_port);
   FA_C_4_0_26 : FA_224 port map( A => q_4_0_26_port, B => q_4_1_26_port, Ci =>
                           q_4_2_26_port, S => q_5_0_26_port, Co => 
                           q_5_1_27_port);
   FA_C_4_0_27 : FA_223 port map( A => q_4_0_27_port, B => q_4_1_27_port, Ci =>
                           q_4_2_27_port, S => q_5_0_27_port, Co => 
                           q_5_1_28_port);
   FA_C_4_0_28 : FA_222 port map( A => q_4_0_28_port, B => q_4_1_28_port, Ci =>
                           q_4_2_28_port, S => q_5_0_28_port, Co => 
                           q_5_1_29_port);
   FA_C_4_0_29 : FA_221 port map( A => q_4_0_29_port, B => q_4_1_29_port, Ci =>
                           q_4_2_29_port, S => q_5_0_29_port, Co => 
                           q_5_1_30_port);
   FA_C_4_0_30 : FA_220 port map( A => q_4_0_30_port, B => q_4_1_30_port, Ci =>
                           q_4_2_30_port, S => q_5_0_30_port, Co => 
                           q_5_1_31_port);
   FA_C_4_0_31 : FA_219 port map( A => q_4_0_31_port, B => q_4_1_31_port, Ci =>
                           q_4_2_31_port, S => q_5_0_31_port, Co => 
                           q_5_1_32_port);
   FA_C_4_0_32 : FA_218 port map( A => q_4_0_32_port, B => q_4_1_32_port, Ci =>
                           q_4_2_32_port, S => q_5_0_32_port, Co => 
                           q_5_1_33_port);
   FA_C_4_0_33 : FA_217 port map( A => q_4_0_33_port, B => q_4_1_33_port, Ci =>
                           q_4_2_33_port, S => q_5_0_33_port, Co => 
                           q_5_1_34_port);
   FA_C_4_0_34 : FA_216 port map( A => q_4_0_34_port, B => q_4_1_34_port, Ci =>
                           q_4_2_34_port, S => q_5_0_34_port, Co => 
                           q_5_1_35_port);
   FA_C_4_0_35 : FA_215 port map( A => q_4_0_35_port, B => q_4_1_35_port, Ci =>
                           q_4_2_35_port, S => q_5_0_35_port, Co => 
                           q_5_1_36_port);
   FA_C_4_0_36 : FA_214 port map( A => q_4_0_36_port, B => q_4_1_36_port, Ci =>
                           q_4_2_36_port, S => q_5_0_36_port, Co => 
                           q_5_1_37_port);
   FA_C_4_0_37 : FA_213 port map( A => q_4_0_37_port, B => q_4_1_37_port, Ci =>
                           q_4_2_37_port, S => q_5_0_37_port, Co => 
                           q_5_1_38_port);
   FA_C_4_0_38 : FA_212 port map( A => q_4_0_38_port, B => q_4_1_38_port, Ci =>
                           q_4_2_38_port, S => q_5_0_38_port, Co_BAR => 
                           q_5_1_39_port);
   FA_C_4_0_39 : FA_211 port map( A => q_4_0_39_port, B => q_4_1_39_port, Ci =>
                           q_4_2_39_port, S => q_5_0_39_port, Co => 
                           q_5_1_40_port);
   FA_C_4_0_40 : FA_210 port map( A => q_4_0_40_port, B => q_4_1_40_port, Ci =>
                           q_4_2_40_port, S => q_5_0_40_port, Co => 
                           q_5_1_41_port);
   FA_C_4_0_41 : FA_209 port map( A => q_4_0_41_port, B => q_4_1_41_port, Ci =>
                           q_4_2_41_port, S => q_5_0_41_port, Co => 
                           q_5_1_42_port);
   FA_C_4_0_42 : FA_208 port map( A => q_4_0_42_port, B => q_4_1_42_port, Ci =>
                           q_4_2_42_port, S => q_5_0_42_port, Co => 
                           q_5_1_43_port);
   FA_C_4_0_43 : FA_207 port map( A => q_4_0_43_port, B => q_4_1_43_port, Ci =>
                           q_4_2_43_port, S => q_5_0_43_port, Co => 
                           q_5_1_44_port);
   FA_C_4_0_44 : FA_206 port map( A => q_4_0_44_port, B => q_4_1_44_port, S => 
                           q_5_0_44_port, Co => q_5_1_45_port, Ci_BAR => 
                           q_4_2_44_port);
   FA_C_4_0_45 : FA_205 port map( A => q_4_0_45_port, B => q_4_1_45_port, S => 
                           q_5_0_45_port, Co => q_5_1_46_port, Ci => 
                           q_4_2_45_port);
   FA_C_4_0_46 : FA_204 port map( A => q_4_0_46_port, B => q_4_1_46_port, S => 
                           q_5_0_46_port, Co => q_5_1_47_port, Ci_BAR => 
                           q_4_2_46_port);
   FA_C_4_0_47 : FA_203 port map( A => q_4_0_47_port, B => q_4_1_47_port, Ci =>
                           q_4_2_47_port, S => q_5_0_47_port, Co => n_2405);
   HA_R_5_0_2 : HA_2 port map( A => q_0_0_2_port, B => q_0_1_2_port, S => 
                           q_6_0_2_port, C => q_6_1_3_port);
   HA_R_5_0_3 : HA_1 port map( A => q_0_0_3_port, B => q_0_1_3_port, S => 
                           q_6_0_3_port, C => q_6_1_4_port);
   FA_C_5_0_4 : FA_188 port map( A => q_5_0_4_port, B => q_0_2_4_port, Ci => 
                           B(5), S => q_6_0_4_port, Co => q_6_1_5_port);
   FA_C_5_0_5 : FA_187 port map( A => q_5_0_5_port, B => q_5_1_5_port, Ci => 
                           q_0_2_5_port, S => q_6_0_5_port, Co => q_6_1_6_port)
                           ;
   FA_C_5_0_6 : FA_186 port map( A => q_5_0_6_port, B => q_5_1_6_port, Ci => 
                           B(7), S => q_6_0_6_port, Co => q_6_1_7_port, clk => 
                           clk);
   FA_C_5_0_7 : FA_185 port map( A => q_5_0_7_port, B => q_5_1_7_port, Ci => 
                           q_0_3_7_port, S => q_6_0_7_port, Co => q_6_1_8_port,
                           clk => clk);
   FA_C_5_0_8 : FA_184 port map( A => q_5_0_8_port, B => q_5_1_8_port, Ci => 
                           B(9), S => q_6_0_8_port, Co => q_6_1_9_port, clk => 
                           clk);
   FA_C_5_0_9 : FA_183 port map( A => q_5_0_9_port, B => q_5_1_9_port, Ci => 
                           q_5_2_9_port, S => q_6_0_9_port, Co => q_6_1_10_port
                           , clk => clk);
   FA_C_5_0_10 : FA_182 port map( A => q_5_0_10_port, B => q_5_1_10_port, Ci =>
                           q_5_2_10_port, S => q_6_0_10_port, Co => 
                           q_6_1_11_port, clk => clk);
   FA_C_5_0_11 : FA_181 port map( A => q_5_0_11_port, B => q_5_1_11_port, Ci =>
                           q_5_2_11_port, S => q_6_0_11_port, Co => 
                           q_6_1_12_port, clk => clk);
   FA_C_5_0_12 : FA_180 port map( A => q_5_0_12_port, B => q_5_1_12_port, Ci =>
                           q_5_2_12_port, S => q_6_0_12_port, Co => 
                           q_6_1_13_port, clk => clk);
   FA_C_5_0_13 : FA_179 port map( A => q_5_0_13_port, B => q_5_1_13_port, Ci =>
                           q_5_2_13_port, S => q_6_0_13_port, Co => 
                           q_6_1_14_port, clk => clk);
   FA_C_5_0_14 : FA_178 port map( A => q_5_0_14_port, B => q_5_1_14_port, Ci =>
                           q_5_2_14_port, S => q_6_0_14_port, Co => 
                           q_6_1_15_port, clk => clk);
   FA_C_5_0_15 : FA_177 port map( A => q_5_0_15_port, B => q_5_1_15_port, Ci =>
                           q_5_2_15_port, S => q_6_0_15_port, Co => 
                           q_6_1_16_port, clk => clk);
   FA_C_5_0_16 : FA_176 port map( A => n193, B => q_5_1_16_port, Ci => 
                           q_5_2_16_port, S => q_6_0_16_port, Co => 
                           q_6_1_17_port);
   FA_C_5_0_17 : FA_175 port map( A => q_5_0_17_port, B => q_5_1_17_port, Ci =>
                           q_5_2_17_port, S => q_6_0_17_port, Co => 
                           q_6_1_18_port);
   FA_C_5_0_18 : FA_174 port map( A => q_5_0_18_port, B => q_5_1_18_port, Ci =>
                           q_5_2_18_port, S => q_6_0_18_port, Co => 
                           q_6_1_19_port);
   FA_C_5_0_19 : FA_173 port map( A => q_5_0_19_port, B => q_5_1_19_port, Ci =>
                           q_5_2_19_port, S => q_6_0_19_port, Co => 
                           q_6_1_20_port);
   FA_C_5_0_20 : FA_172 port map( A => q_5_0_20_port, B => q_5_1_20_port, Ci =>
                           q_5_2_20_port, S => q_6_0_20_port, Co => 
                           q_6_1_21_port);
   FA_C_5_0_21 : FA_171 port map( A => q_5_0_21_port, B => q_5_1_21_port, Ci =>
                           q_5_2_21_port, S => q_6_0_21_port, Co => 
                           q_6_1_22_port);
   FA_C_5_0_22 : FA_170 port map( A => q_5_0_22_port, B => q_5_1_22_port, Ci =>
                           q_5_2_22_port, S => q_6_0_22_port, Co => 
                           q_6_1_23_port);
   FA_C_5_0_23 : FA_169 port map( A => q_5_0_23_port, B => q_5_1_23_port, Ci =>
                           q_5_2_23_port, S => q_6_0_23_port, Co => 
                           q_6_1_24_port);
   FA_C_5_0_24 : FA_168 port map( A => q_5_0_24_port, B => q_5_1_24_port, Ci =>
                           q_5_2_24_port, S => q_6_0_24_port, Co => 
                           q_6_1_25_port);
   FA_C_5_0_25 : FA_167 port map( A => q_5_0_25_port, B => q_5_1_25_port, Ci =>
                           q_5_2_25_port, S => q_6_0_25_port, Co => 
                           q_6_1_26_port);
   FA_C_5_0_26 : FA_166 port map( A => q_5_0_26_port, B => q_5_1_26_port, Ci =>
                           q_5_2_26_port, S => q_6_0_26_port, Co => n177);
   FA_C_5_0_27 : FA_165 port map( A => q_5_0_27_port, B => q_5_1_27_port, Ci =>
                           q_5_2_27_port, S => q_6_0_27_port, Co => 
                           q_6_1_28_port);
   FA_C_5_0_28 : FA_164 port map( A => q_5_0_28_port, B => q_5_1_28_port, Ci =>
                           q_5_2_28_port, S => q_6_0_28_port, Co => n175);
   FA_C_5_0_29 : FA_163 port map( A => q_5_0_29_port, B => q_5_1_29_port, Ci =>
                           q_5_2_29_port, S => q_6_0_29_port, Co => 
                           q_6_1_30_port);
   FA_C_5_0_30 : FA_162 port map( A => q_5_0_30_port, B => q_5_1_30_port, Ci =>
                           q_5_2_30_port, S => q_6_0_30_port, Co => 
                           q_6_1_31_port);
   FA_C_5_0_31 : FA_161 port map( A => q_5_0_31_port, B => q_5_1_31_port, Ci =>
                           q_5_2_31_port, S => q_6_0_31_port, Co => 
                           q_6_1_32_port);
   FA_C_5_0_32 : FA_160 port map( A => q_5_0_32_port, B => q_5_1_32_port, Ci =>
                           q_5_2_32_port, S => q_6_0_32_port, Co => n173);
   FA_C_5_0_33 : FA_159 port map( A => q_5_0_33_port, B => q_5_1_33_port, Ci =>
                           q_5_2_33_port, S => n178, Co => q_6_1_34_port);
   FA_C_5_0_34 : FA_158 port map( A => q_5_0_34_port, B => q_5_1_34_port, Ci =>
                           q_5_2_34_port, S => q_6_0_34_port, Co => n174);
   FA_C_5_0_35 : FA_157 port map( A => q_5_0_35_port, B => q_5_1_35_port, Ci =>
                           net102732, S => q_6_0_35_port, Co => q_6_1_36_port);
   FA_C_5_0_36 : FA_156 port map( A => q_5_0_36_port, B => q_5_1_36_port, Ci =>
                           net102731, S => q_6_0_36_port, Co => q_6_1_37_port);
   FA_C_5_0_37 : FA_155 port map( A => q_5_0_37_port, B => q_5_1_37_port, Ci =>
                           net102730, S => q_6_0_37_port, Co => q_6_1_38_port);
   FA_C_5_0_38 : FA_154 port map( A => q_5_0_38_port, B => q_5_1_38_port, Ci =>
                           net102729, S => q_6_0_38_port, Co => q_6_1_39_port);
   FA_C_5_0_39 : FA_153 port map( A => q_5_0_39_port, Ci => net102728, S => 
                           n176, Co => q_6_1_40_port, B_BAR => q_5_1_39_port);
   FA_C_5_0_40 : FA_152 port map( A => q_5_0_40_port, B => q_5_1_40_port, Ci =>
                           net102727, S => q_6_0_40_port, Co => q_6_1_41_port);
   FA_C_5_0_41 : FA_151 port map( A => q_5_0_41_port, B => q_5_1_41_port, Ci =>
                           net102726, S => q_6_0_41_port, Co => q_6_1_42_port);
   FA_C_5_0_42 : FA_150 port map( A => q_5_0_42_port, B => q_5_1_42_port, Ci =>
                           net102725, S => q_6_0_42_port, Co => q_6_1_43_port);
   FA_C_5_0_43 : FA_149 port map( A => q_5_0_43_port, B => q_5_1_43_port, Ci =>
                           q_5_2_43_port, S => q_6_0_43_port, Co => 
                           q_6_1_44_port);
   FA_C_5_0_44 : FA_148 port map( A => q_5_0_44_port, B => q_5_1_44_port, Ci =>
                           q_5_2_44_port, S => q_6_0_44_port, Co => 
                           q_6_1_45_port);
   FA_C_5_0_45 : FA_147 port map( A => q_5_0_45_port, B => q_5_1_45_port, Ci =>
                           q_5_2_45_port, S => q_6_0_45_port, Co => 
                           q_6_1_46_port);
   FA_C_5_0_46 : FA_146 port map( A => q_5_0_46_port, B => q_5_1_46_port, Ci =>
                           net102724, S => q_6_0_46_port, Co => q_6_1_47_port);
   FA_C_5_0_47 : FA_145 port map( A => q_5_0_47_port, B => q_5_1_47_port, Ci =>
                           q_5_2_47_port, S => q_6_0_47_port, Co => n_2406);
   P4_ADDER_0 : P4_ADDER_NBIT64_NBIT_PER_BLOCK2_NBLOCKS32 port map( A(63) => 
                           n140, A(62) => n141, A(61) => n142, A(60) => n143, 
                           A(59) => n144, A(58) => n145, A(57) => n146, A(56) 
                           => n147, A(55) => n148, A(54) => n149, A(53) => n150
                           , A(52) => n151, A(51) => n152, A(50) => n153, A(49)
                           => n154, A(48) => n155, A(47) => q_6_0_47_port, 
                           A(46) => q_6_0_46_port, A(45) => q_6_0_45_port, 
                           A(44) => q_6_0_44_port, A(43) => q_6_0_43_port, 
                           A(42) => q_6_0_42_port, A(41) => q_6_0_41_port, 
                           A(40) => q_6_0_40_port, A(39) => n176, A(38) => 
                           q_6_0_38_port, A(37) => q_6_0_37_port, A(36) => 
                           q_6_0_36_port, A(35) => q_6_0_35_port, A(34) => 
                           q_6_0_34_port, A(33) => n178, A(32) => q_6_0_32_port
                           , A(31) => q_6_0_31_port, A(30) => q_6_0_30_port, 
                           A(29) => q_6_0_29_port, A(28) => q_6_0_28_port, 
                           A(27) => q_6_0_27_port, A(26) => q_6_0_26_port, 
                           A(25) => q_6_0_25_port, A(24) => q_6_0_24_port, 
                           A(23) => q_6_0_23_port, A(22) => q_6_0_22_port, 
                           A(21) => q_6_0_21_port, A(20) => q_6_0_20_port, 
                           A(19) => q_6_0_19_port, A(18) => q_6_0_18_port, 
                           A(17) => q_6_0_17_port, A(16) => q_6_0_16_port, 
                           A(15) => q_6_0_15_port, A(14) => q_6_0_14_port, 
                           A(13) => q_6_0_13_port, A(12) => q_6_0_12_port, 
                           A(11) => q_6_0_11_port, A(10) => q_6_0_10_port, A(9)
                           => q_6_0_9_port, A(8) => q_6_0_8_port, A(7) => 
                           q_6_0_7_port, A(6) => q_6_0_6_port, A(5) => 
                           q_6_0_5_port, A(4) => q_6_0_4_port, A(3) => 
                           q_6_0_3_port, A(2) => q_6_0_2_port, A(1) => 
                           q_0_0_1_port, A(0) => q_0_0_0_port, B(63) => n156, 
                           B(62) => n157, B(61) => n158, B(60) => n159, B(59) 
                           => n160, B(58) => n161, B(57) => n162, B(56) => n163
                           , B(55) => n164, B(54) => n165, B(53) => n166, B(52)
                           => n167, B(51) => n168, B(50) => n169, B(49) => n170
                           , B(48) => n171, B(47) => q_6_1_47_port, B(46) => 
                           q_6_1_46_port, B(45) => q_6_1_45_port, B(44) => 
                           q_6_1_44_port, B(43) => q_6_1_43_port, B(42) => 
                           q_6_1_42_port, B(41) => q_6_1_41_port, B(40) => 
                           q_6_1_40_port, B(39) => q_6_1_39_port, B(38) => 
                           q_6_1_38_port, B(37) => q_6_1_37_port, B(36) => 
                           q_6_1_36_port, B(35) => n174, B(34) => q_6_1_34_port
                           , B(33) => n173, B(32) => q_6_1_32_port, B(31) => 
                           q_6_1_31_port, B(30) => q_6_1_30_port, B(29) => n175
                           , B(28) => q_6_1_28_port, B(27) => n177, B(26) => 
                           q_6_1_26_port, B(25) => q_6_1_25_port, B(24) => 
                           q_6_1_24_port, B(23) => q_6_1_23_port, B(22) => 
                           q_6_1_22_port, B(21) => q_6_1_21_port, B(20) => 
                           q_6_1_20_port, B(19) => q_6_1_19_port, B(18) => 
                           q_6_1_18_port, B(17) => q_6_1_17_port, B(16) => 
                           q_6_1_16_port, B(15) => q_6_1_15_port, B(14) => 
                           q_6_1_14_port, B(13) => q_6_1_13_port, B(12) => 
                           q_6_1_12_port, B(11) => q_6_1_11_port, B(10) => 
                           q_6_1_10_port, B(9) => q_6_1_9_port, B(8) => 
                           q_6_1_8_port, B(7) => q_6_1_7_port, B(6) => 
                           q_6_1_6_port, B(5) => q_6_1_5_port, B(4) => 
                           q_6_1_4_port, B(3) => q_6_1_3_port, B(2) => B(3), 
                           B(1) => X_Logic0_port, B(0) => B(1), Cin => 
                           X_Logic0_port, S(63) => n_2407, S(62) => n_2408, 
                           S(61) => n_2409, S(60) => n_2410, S(59) => n_2411, 
                           S(58) => n_2412, S(57) => n_2413, S(56) => n_2414, 
                           S(55) => n_2415, S(54) => n_2416, S(53) => n_2417, 
                           S(52) => n_2418, S(51) => n_2419, S(50) => n_2420, 
                           S(49) => n_2421, S(48) => n_2422, S(47) => C(47), 
                           S(46) => C(46), S(45) => C(45), S(44) => C(44), 
                           S(43) => C(43), S(42) => C(42), S(41) => C(41), 
                           S(40) => C(40), S(39) => C(39), S(38) => C(38), 
                           S(37) => C(37), S(36) => C(36), S(35) => C(35), 
                           S(34) => C(34), S(33) => C(33), S(32) => C(32), 
                           S(31) => C(31), S(30) => C(30), S(29) => C(29), 
                           S(28) => C(28), S(27) => C(27), S(26) => C(26), 
                           S(25) => C(25), S(24) => C(24), S(23) => C(23), 
                           S(22) => C(22), S(21) => n_2423, S(20) => n_2424, 
                           S(19) => n_2425, S(18) => n_2426, S(17) => n_2427, 
                           S(16) => n_2428, S(15) => n_2429, S(14) => n_2430, 
                           S(13) => n_2431, S(12) => n_2432, S(11) => n_2433, 
                           S(10) => n_2434, S(9) => n_2435, S(8) => n_2436, 
                           S(7) => n_2437, S(6) => n_2438, S(5) => n_2439, S(4)
                           => n_2440, S(3) => n_2441, S(2) => n_2442, S(1) => 
                           n_2443, S(0) => n_2444, Cout => n_2445, clk => clk);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity UnpackFP_1 is

   port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector 
         (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, isNaN,
         isINF, isZ, isDN : out std_logic);

end UnpackFP_1;

architecture SYN_UnpackFP of UnpackFP_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N13, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13_port, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n_2446, n_2447, n_2448, 
      n_2449, n_2450, n_2451, n_2452, n_2453 : std_logic;

begin
   SIG <= ( n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, N13
      , FP(22), FP(21), FP(20), FP(19), FP(18), FP(17), FP(16), FP(15), FP(14),
      FP(13), FP(12), FP(11), FP(10), FP(9), FP(8), FP(7), FP(6), FP(5), FP(4),
      FP(3), FP(2), FP(1), FP(0) );
   EXP <= ( FP(30), FP(29), FP(28), FP(27), FP(26), FP(25), FP(24), FP(23) );
   SIGN <= FP(31);
   
   U2 : NAND4_X1 port map( A1 => n24, A2 => n23, A3 => n22, A4 => n21, ZN => 
                           n35);
   U3 : NOR2_X1 port map( A1 => FP(0), A2 => FP(1), ZN => n24);
   U4 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => n22);
   U5 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U6 : NOR2_X1 port map( A1 => FP(10), A2 => FP(9), ZN => n3);
   U7 : INV_X1 port map( A => FP(19), ZN => n17);
   U8 : INV_X1 port map( A => FP(20), ZN => n16);
   U9 : NOR2_X1 port map( A1 => FP(18), A2 => FP(17), ZN => n18);
   U10 : INV_X1 port map( A => FP(13), ZN => n12);
   U11 : INV_X1 port map( A => FP(14), ZN => n11);
   U12 : NOR2_X1 port map( A1 => FP(12), A2 => FP(11), ZN => n13_port);
   U13 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n23);
   U14 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n9);
   U15 : NAND4_X1 port map( A1 => n6, A2 => n5, A3 => n4, A4 => n3, ZN => n10);
   U16 : INV_X1 port map( A => FP(4), ZN => n7);
   U17 : NOR2_X1 port map( A1 => FP(3), A2 => FP(2), ZN => n8);
   U18 : NOR2_X1 port map( A1 => FP(5), A2 => FP(6), ZN => n6);
   U19 : OR2_X1 port map( A1 => FP(22), A2 => FP(21), ZN => n19);
   U20 : OR2_X1 port map( A1 => FP(16), A2 => FP(15), ZN => n14);
   U21 : INV_X1 port map( A => FP(8), ZN => n4);
   U22 : INV_X1 port map( A => FP(7), ZN => n5);
   U23 : NOR4_X1 port map( A1 => FP(27), A2 => FP(28), A3 => FP(29), A4 => 
                           FP(30), ZN => n2);
   U24 : NOR4_X1 port map( A1 => FP(23), A2 => FP(24), A3 => FP(25), A4 => 
                           FP(26), ZN => n1);
   U25 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => N13);
   U26 : NAND3_X1 port map( A1 => n13_port, A2 => n12, A3 => n11, ZN => n15);
   U27 : NAND3_X1 port map( A1 => n18, A2 => n17, A3 => n16, ZN => n20);
   U28 : INV_X1 port map( A => n35, ZN => n37);
   U30 : NOR2_X1 port map( A1 => N13, A2 => n35, ZN => isZ);
   U31 : INV_X1 port map( A => FP(28), ZN => n28);
   U32 : INV_X1 port map( A => FP(27), ZN => n27);
   U33 : INV_X1 port map( A => FP(30), ZN => n26);
   U34 : INV_X1 port map( A => FP(29), ZN => n25);
   U35 : NOR4_X1 port map( A1 => n28, A2 => n27, A3 => n26, A4 => n25, ZN => 
                           n34);
   U36 : INV_X1 port map( A => FP(24), ZN => n32);
   U37 : INV_X1 port map( A => FP(23), ZN => n31);
   U38 : INV_X1 port map( A => FP(26), ZN => n30);
   U39 : INV_X1 port map( A => FP(25), ZN => n29);
   U40 : NOR4_X1 port map( A1 => n32, A2 => n31, A3 => n30, A4 => n29, ZN => 
                           n33);
   U41 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => n36);
   U42 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => isINF);
   U43 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => isNaN);

end SYN_UnpackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity UnpackFP_0 is

   port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector 
         (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, isNaN,
         isINF, isZ, isDN : out std_logic);

end UnpackFP_0;

architecture SYN_UnpackFP of UnpackFP_0 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N13, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13_port, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n_2455, n_2456, n_2457, 
      n_2458, n_2459, n_2460, n_2461, n_2462 : std_logic;

begin
   SIG <= ( n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, N13
      , FP(22), FP(21), FP(20), FP(19), FP(18), FP(17), FP(16), FP(15), FP(14),
      FP(13), FP(12), FP(11), FP(10), FP(9), FP(8), FP(7), FP(6), FP(5), FP(4),
      FP(3), FP(2), FP(1), FP(0) );
   EXP <= ( FP(30), FP(29), FP(28), FP(27), FP(26), FP(25), FP(24), FP(23) );
   SIGN <= FP(31);
   
   U2 : NAND4_X1 port map( A1 => n24, A2 => n23, A3 => n22, A4 => n21, ZN => 
                           n35);
   U3 : NOR2_X1 port map( A1 => FP(0), A2 => FP(1), ZN => n24);
   U4 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => n22);
   U5 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U6 : NOR2_X1 port map( A1 => FP(10), A2 => FP(9), ZN => n3);
   U7 : INV_X1 port map( A => FP(19), ZN => n17);
   U8 : INV_X1 port map( A => FP(20), ZN => n16);
   U9 : NOR2_X1 port map( A1 => FP(18), A2 => FP(17), ZN => n18);
   U10 : INV_X1 port map( A => FP(13), ZN => n12);
   U11 : INV_X1 port map( A => FP(14), ZN => n11);
   U12 : NOR2_X1 port map( A1 => FP(12), A2 => FP(11), ZN => n13_port);
   U13 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n23);
   U14 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n9);
   U15 : NAND4_X1 port map( A1 => n6, A2 => n5, A3 => n4, A4 => n3, ZN => n10);
   U16 : INV_X1 port map( A => FP(4), ZN => n7);
   U17 : NOR2_X1 port map( A1 => FP(3), A2 => FP(2), ZN => n8);
   U18 : NOR2_X1 port map( A1 => FP(5), A2 => FP(6), ZN => n6);
   U19 : OR2_X1 port map( A1 => FP(22), A2 => FP(21), ZN => n19);
   U20 : OR2_X1 port map( A1 => FP(16), A2 => FP(15), ZN => n14);
   U21 : INV_X1 port map( A => FP(8), ZN => n4);
   U22 : INV_X1 port map( A => FP(7), ZN => n5);
   U23 : NOR4_X1 port map( A1 => FP(27), A2 => FP(28), A3 => FP(29), A4 => 
                           FP(30), ZN => n2);
   U24 : NOR4_X1 port map( A1 => FP(23), A2 => FP(24), A3 => FP(25), A4 => 
                           FP(26), ZN => n1);
   U26 : NAND3_X1 port map( A1 => n13_port, A2 => n12, A3 => n11, ZN => n15);
   U27 : NAND3_X1 port map( A1 => n18, A2 => n17, A3 => n16, ZN => n20);
   U28 : INV_X1 port map( A => n35, ZN => n37);
   U30 : NOR2_X1 port map( A1 => N13, A2 => n35, ZN => isZ);
   U31 : INV_X1 port map( A => FP(28), ZN => n28);
   U32 : INV_X1 port map( A => FP(27), ZN => n27);
   U33 : INV_X1 port map( A => FP(30), ZN => n26);
   U34 : INV_X1 port map( A => FP(29), ZN => n25);
   U35 : NOR4_X1 port map( A1 => n28, A2 => n27, A3 => n26, A4 => n25, ZN => 
                           n34);
   U36 : INV_X1 port map( A => FP(24), ZN => n32);
   U37 : INV_X1 port map( A => FP(23), ZN => n31);
   U38 : INV_X1 port map( A => FP(26), ZN => n30);
   U39 : INV_X1 port map( A => FP(25), ZN => n29);
   U40 : NOR4_X1 port map( A1 => n32, A2 => n31, A3 => n30, A4 => n29, ZN => 
                           n33);
   U41 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => n36);
   U42 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => isINF);
   U43 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => isNaN);
   U25 : NAND2_X2 port map( A1 => n2, A2 => n1, ZN => N13);

end SYN_UnpackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage4 is

   port( EXP_neg : in std_logic;  EXP_out_round : in std_logic_vector (7 downto
         0);  EXP_pos, SIGN_out : in std_logic;  SIG_out_round : in 
         std_logic_vector (27 downto 0);  clk, isINF_tab, isNaN, isZ_tab : in 
         std_logic;  FP_Z : out std_logic_vector (31 downto 0));

end FPmul_stage4;

architecture SYN_struct of FPmul_stage4 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component PackFP
      port( SIGN : in std_logic;  EXP : in std_logic_vector (7 downto 0);  SIG 
            : in std_logic_vector (22 downto 0);  isNaN, isINF, isZ : in 
            std_logic;  FP : out std_logic_vector (31 downto 0);  clk : in 
            std_logic);
   end component;
   
   component FPnormalize_SIG_width28_1
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
            std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n171, SIG_out_norm2_26_port, SIG_out_22_port, SIG_out_21_port, 
      SIG_out_20_port, SIG_out_19_port, SIG_out_18_port, SIG_out_17_port, 
      SIG_out_16_port, SIG_out_15_port, SIG_out_14_port, SIG_out_13_port, 
      SIG_out_12_port, SIG_out_11_port, SIG_out_10_port, SIG_out_9_port, 
      SIG_out_8_port, SIG_out_7_port, SIG_out_6_port, SIG_out_5_port, 
      SIG_out_4_port, SIG_out_3_port, SIG_out_2_port, SIG_out_1_port, 
      SIG_out_0_port, EXP_out_7_port, EXP_out_6_port, EXP_out_5_port, 
      EXP_out_4_port, EXP_out_3_port, EXP_out_2_port, EXP_out_1_port, 
      EXP_out_0_port, isINF, n1, n5, n9, n13, n17, n18, n19, n20, n21, n26, n28
      , n29, n30, n31, n32, n33, n69, n70, n71, n72, n74, n75, n76, n77, n78, 
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, n97, n98, n99, n100, n101, n102, n168, n169, n170, n174,
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n_2467, n_2468, n_2469, n_2470, n_2471, 
      n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, 
      n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, 
      n_2490, n_2491, n_2492, n_2493 : std_logic;

begin
   
   U9 : INV_X1 port map( A => isINF_tab, ZN => n31);
   U10 : INV_X1 port map( A => EXP_pos, ZN => n29);
   U15 : NOR3_X1 port map( A1 => n79, A2 => n80, A3 => n81, ZN => n1);
   U16 : NAND4_X1 port map( A1 => n185, A2 => n184, A3 => n177, A4 => n1, ZN =>
                           n20);
   U20 : NOR3_X1 port map( A1 => n85, A2 => n86, A3 => n87, ZN => n5);
   U21 : NAND4_X1 port map( A1 => n176, A2 => n186, A3 => n187, A4 => n5, ZN =>
                           n19);
   U25 : NOR3_X1 port map( A1 => n91, A2 => n92, A3 => n93, ZN => n9);
   U26 : NAND4_X1 port map( A1 => n182, A2 => n174, A3 => n175, A4 => n9, ZN =>
                           n18);
   U30 : NOR3_X1 port map( A1 => n100, A2 => n101, A3 => n102, ZN => n13);
   U31 : NAND4_X1 port map( A1 => n178, A2 => n180, A3 => n183, A4 => n13, ZN 
                           => n17);
   U32 : NOR4_X1 port map( A1 => n20, A2 => n19, A3 => n18, A4 => n17, ZN => 
                           n21);
   U34 : INV_X1 port map( A => n30, ZN => n33);
   MY_CLK_r_REG242_S4 : DFF_X1 port map( D => n74, CK => clk, Q => n_2467, QN 
                           => n179);
   n168 <= '0';
   n169 <= '0';
   n170 <= '0';
   U3 : AND2_X1 port map( A1 => EXP_out_2_port, A2 => n77, ZN => n26);
   U4 : OR2_X1 port map( A1 => n21, A2 => n69, ZN => n191);
   U5 : AND2_X1 port map( A1 => n26, A2 => n78, ZN => n181);
   U6 : AND2_X1 port map( A1 => EXP_out_3_port, A2 => EXP_out_4_port, ZN => 
                           n188);
   U7 : NAND4_X1 port map( A1 => n188, A2 => EXP_out_6_port, A3 => 
                           EXP_out_5_port, A4 => n181, ZN => n28);
   U8 : NAND2_X1 port map( A1 => n190, A2 => n189, ZN => n32);
   U11 : OR2_X1 port map( A1 => EXP_out_7_port, A2 => n179, ZN => n189);
   U12 : NAND2_X1 port map( A1 => n28, A2 => EXP_out_7_port, ZN => n190);
   U13 : AOI21_X1 port map( B1 => n32, B2 => n75, A => n33, ZN => isINF);
   U14 : AOI21_X1 port map( B1 => EXP_out_7_port, B2 => n71, A => n191, ZN => 
                           n30);
   I1 : FPnormalize_SIG_width28_1 port map( SIG_in(27) => SIG_out_round(27), 
                           SIG_in(26) => SIG_out_round(26), SIG_in(25) => 
                           SIG_out_round(25), SIG_in(24) => SIG_out_round(24), 
                           SIG_in(23) => SIG_out_round(23), SIG_in(22) => 
                           SIG_out_round(22), SIG_in(21) => SIG_out_round(21), 
                           SIG_in(20) => SIG_out_round(20), SIG_in(19) => 
                           SIG_out_round(19), SIG_in(18) => SIG_out_round(18), 
                           SIG_in(17) => SIG_out_round(17), SIG_in(16) => 
                           SIG_out_round(16), SIG_in(15) => SIG_out_round(15), 
                           SIG_in(14) => SIG_out_round(14), SIG_in(13) => 
                           SIG_out_round(13), SIG_in(12) => SIG_out_round(12), 
                           SIG_in(11) => SIG_out_round(11), SIG_in(10) => 
                           SIG_out_round(10), SIG_in(9) => SIG_out_round(9), 
                           SIG_in(8) => SIG_out_round(8), SIG_in(7) => 
                           SIG_out_round(7), SIG_in(6) => SIG_out_round(6), 
                           SIG_in(5) => SIG_out_round(5), SIG_in(4) => 
                           SIG_out_round(4), SIG_in(3) => SIG_out_round(3), 
                           SIG_in(2) => n168, SIG_in(1) => n169, SIG_in(0) => 
                           n170, EXP_in(7) => EXP_out_round(7), EXP_in(6) => 
                           EXP_out_round(6), EXP_in(5) => EXP_out_round(5), 
                           EXP_in(4) => EXP_out_round(4), EXP_in(3) => 
                           EXP_out_round(3), EXP_in(2) => EXP_out_round(2), 
                           EXP_in(1) => EXP_out_round(1), EXP_in(0) => 
                           EXP_out_round(0), SIG_out(27) => n_2468, SIG_out(26)
                           => SIG_out_norm2_26_port, SIG_out(25) => 
                           SIG_out_22_port, SIG_out(24) => SIG_out_21_port, 
                           SIG_out(23) => SIG_out_20_port, SIG_out(22) => 
                           SIG_out_19_port, SIG_out(21) => SIG_out_18_port, 
                           SIG_out(20) => SIG_out_17_port, SIG_out(19) => 
                           SIG_out_16_port, SIG_out(18) => SIG_out_15_port, 
                           SIG_out(17) => SIG_out_14_port, SIG_out(16) => 
                           SIG_out_13_port, SIG_out(15) => SIG_out_12_port, 
                           SIG_out(14) => SIG_out_11_port, SIG_out(13) => 
                           SIG_out_10_port, SIG_out(12) => SIG_out_9_port, 
                           SIG_out(11) => SIG_out_8_port, SIG_out(10) => 
                           SIG_out_7_port, SIG_out(9) => SIG_out_6_port, 
                           SIG_out(8) => SIG_out_5_port, SIG_out(7) => 
                           SIG_out_4_port, SIG_out(6) => SIG_out_3_port, 
                           SIG_out(5) => SIG_out_2_port, SIG_out(4) => 
                           SIG_out_1_port, SIG_out(3) => SIG_out_0_port, 
                           SIG_out(2) => n_2469, SIG_out(1) => n_2470, 
                           SIG_out(0) => n_2471, EXP_out(7) => EXP_out_7_port, 
                           EXP_out(6) => EXP_out_6_port, EXP_out(5) => 
                           EXP_out_5_port, EXP_out(4) => EXP_out_4_port, 
                           EXP_out(3) => EXP_out_3_port, EXP_out(2) => 
                           EXP_out_2_port, EXP_out(1) => EXP_out_1_port, 
                           EXP_out(0) => EXP_out_0_port, clk => clk);
   I3 : PackFP port map( SIGN => SIGN_out, EXP(7) => EXP_out_7_port, EXP(6) => 
                           EXP_out_6_port, EXP(5) => EXP_out_5_port, EXP(4) => 
                           EXP_out_4_port, EXP(3) => EXP_out_3_port, EXP(2) => 
                           EXP_out_2_port, EXP(1) => n78, EXP(0) => n77, 
                           SIG(22) => n101, SIG(21) => n100, SIG(20) => n99, 
                           SIG(19) => n98, SIG(18) => n97, SIG(17) => n96, 
                           SIG(16) => n95, SIG(15) => n94, SIG(14) => n93, 
                           SIG(13) => n92, SIG(12) => n91, SIG(11) => n90, 
                           SIG(10) => n89, SIG(9) => n88, SIG(8) => n87, SIG(7)
                           => n86, SIG(6) => n85, SIG(5) => n84, SIG(4) => n83,
                           SIG(3) => n82, SIG(2) => n81, SIG(1) => n80, SIG(0) 
                           => n79, isNaN => isNaN, isINF => isINF, isZ => n33, 
                           FP(31) => n171, FP(30) => FP_Z(30), FP(29) => 
                           FP_Z(29), FP(28) => FP_Z(28), FP(27) => FP_Z(27), 
                           FP(26) => FP_Z(26), FP(25) => FP_Z(25), FP(24) => 
                           FP_Z(24), FP(23) => FP_Z(23), FP(22) => FP_Z(22), 
                           FP(21) => FP_Z(21), FP(20) => FP_Z(20), FP(19) => 
                           FP_Z(19), FP(18) => FP_Z(18), FP(17) => FP_Z(17), 
                           FP(16) => FP_Z(16), FP(15) => FP_Z(15), FP(14) => 
                           FP_Z(14), FP(13) => FP_Z(13), FP(12) => FP_Z(12), 
                           FP(11) => FP_Z(11), FP(10) => FP_Z(10), FP(9) => 
                           FP_Z(9), FP(8) => FP_Z(8), FP(7) => FP_Z(7), FP(6) 
                           => FP_Z(6), FP(5) => FP_Z(5), FP(4) => FP_Z(4), 
                           FP(3) => FP_Z(3), FP(2) => FP_Z(2), FP(1) => FP_Z(1)
                           , FP(0) => FP_Z(0), clk => clk);
   MY_CLK_r_REG47_S4 : DFF_X1 port map( D => SIG_out_10_port, CK => clk, Q => 
                           n89, QN => n186);
   MY_CLK_r_REG46_S4 : DFF_X1 port map( D => SIG_out_11_port, CK => clk, Q => 
                           n90, QN => n176);
   MY_CLK_r_REG42_S4 : DFF_X1 port map( D => SIG_out_15_port, CK => clk, Q => 
                           n94, QN => n175);
   MY_CLK_r_REG41_S4 : DFF_X1 port map( D => SIG_out_16_port, CK => clk, Q => 
                           n95, QN => n174);
   MY_CLK_r_REG40_S4 : DFF_X1 port map( D => SIG_out_17_port, CK => clk, Q => 
                           n96, QN => n182);
   MY_CLK_r_REG39_S4 : DFF_X1 port map( D => SIG_out_18_port, CK => clk, Q => 
                           n97, QN => n183);
   MY_CLK_r_REG38_S4 : DFF_X1 port map( D => SIG_out_19_port, CK => clk, Q => 
                           n98, QN => n180);
   MY_CLK_r_REG37_S4 : DFF_X1 port map( D => SIG_out_20_port, CK => clk, Q => 
                           n99, QN => n178);
   MY_CLK_r_REG31_S4 : DFF_X1 port map( D => SIG_out_3_port, CK => clk, Q => 
                           n82, QN => n177);
   MY_CLK_r_REG30_S4 : DFF_X1 port map( D => SIG_out_4_port, CK => clk, Q => 
                           n83, QN => n184);
   MY_CLK_r_REG29_S4 : DFF_X1 port map( D => SIG_out_5_port, CK => clk, Q => 
                           n84, QN => n185);
   MY_CLK_r_REG25_S4 : DFF_X1 port map( D => SIG_out_9_port, CK => clk, Q => 
                           n88, QN => n187);
   MY_CLK_r_REG241_S3 : DFF_X1 port map( D => n29, CK => clk, Q => n74, QN => 
                           n_2472);
   MY_CLK_r_REG239_S4 : DFF_X1 port map( D => n72, CK => clk, Q => n71, QN => 
                           n_2473);
   MY_CLK_r_REG238_S3 : DFF_X1 port map( D => EXP_neg, CK => clk, Q => n72, QN 
                           => n_2474);
   MY_CLK_r_REG45_S4 : DFF_X1 port map( D => SIG_out_12_port, CK => clk, Q => 
                           n91, QN => n_2475);
   MY_CLK_r_REG44_S4 : DFF_X1 port map( D => SIG_out_13_port, CK => clk, Q => 
                           n92, QN => n_2476);
   MY_CLK_r_REG43_S4 : DFF_X1 port map( D => SIG_out_14_port, CK => clk, Q => 
                           n93, QN => n_2477);
   MY_CLK_r_REG36_S4 : DFF_X1 port map( D => SIG_out_21_port, CK => clk, Q => 
                           n100, QN => n_2478);
   MY_CLK_r_REG35_S4 : DFF_X1 port map( D => EXP_out_0_port, CK => clk, Q => 
                           n77, QN => n_2479);
   MY_CLK_r_REG34_S4 : DFF_X1 port map( D => SIG_out_0_port, CK => clk, Q => 
                           n79, QN => n_2480);
   MY_CLK_r_REG33_S4 : DFF_X1 port map( D => SIG_out_1_port, CK => clk, Q => 
                           n80, QN => n_2481);
   MY_CLK_r_REG32_S4 : DFF_X1 port map( D => SIG_out_2_port, CK => clk, Q => 
                           n81, QN => n_2482);
   MY_CLK_r_REG28_S4 : DFF_X1 port map( D => SIG_out_6_port, CK => clk, Q => 
                           n85, QN => n_2483);
   MY_CLK_r_REG27_S4 : DFF_X1 port map( D => SIG_out_7_port, CK => clk, Q => 
                           n86, QN => n_2484);
   MY_CLK_r_REG26_S4 : DFF_X1 port map( D => SIG_out_8_port, CK => clk, Q => 
                           n87, QN => n_2485);
   MY_CLK_r_REG24_S4 : DFF_X1 port map( D => SIG_out_22_port, CK => clk, Q => 
                           n101, QN => n_2486);
   MY_CLK_r_REG23_S4 : DFF_X1 port map( D => SIG_out_norm2_26_port, CK => clk, 
                           Q => n102, QN => n_2487);
   MY_CLK_r_REG19_S4 : DFF_X1 port map( D => EXP_out_1_port, CK => clk, Q => 
                           n78, QN => n_2488);
   MY_CLK_r_REG15_S4 : DFF_X1 port map( D => n76, CK => clk, Q => n75, QN => 
                           n_2489);
   MY_CLK_r_REG14_S3 : DFF_X1 port map( D => n31, CK => clk, Q => n76, QN => 
                           n_2490);
   MY_CLK_r_REG11_S4 : DFF_X1 port map( D => n70, CK => clk, Q => n69, QN => 
                           n_2491);
   MY_CLK_r_REG10_S3 : DFF_X1 port map( D => isZ_tab, CK => clk, Q => n70, QN 
                           => n_2492);
   MY_CLK_r_REG2_S3 : DFF_X1 port map( D => n171, CK => clk, Q => FP_Z(31), QN 
                           => n_2493);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage3 is

   port( EXP_in : in std_logic_vector (7 downto 0);  EXP_neg_stage2, 
         EXP_pos_stage2, SIGN_out_stage2 : in std_logic;  SIG_in : in 
         std_logic_vector (27 downto 0);  clk, isINF_stage2, isNaN_stage2, 
         isZ_tab_stage2 : in std_logic;  EXP_neg : out std_logic;  
         EXP_out_round : out std_logic_vector (7 downto 0);  EXP_pos, SIGN_out 
         : out std_logic;  SIG_out_round : out std_logic_vector (27 downto 0); 
         isINF_tab, isNaN, isZ_tab : out std_logic);

end FPmul_stage3;

architecture SYN_struct of FPmul_stage3 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FPround_SIG_width28
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
            std_logic);
   end component;
   
   component FPnormalize_SIG_width28_0
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
            std_logic);
   end component;
   
   signal SIG_out_norm_27_port, SIG_out_norm_26_port, SIG_out_norm_25_port, 
      SIG_out_norm_24_port, SIG_out_norm_23_port, SIG_out_norm_22_port, 
      SIG_out_norm_21_port, SIG_out_norm_20_port, SIG_out_norm_19_port, 
      SIG_out_norm_18_port, SIG_out_norm_17_port, SIG_out_norm_16_port, 
      SIG_out_norm_15_port, SIG_out_norm_14_port, SIG_out_norm_13_port, 
      SIG_out_norm_12_port, SIG_out_norm_11_port, SIG_out_norm_10_port, 
      SIG_out_norm_9_port, SIG_out_norm_8_port, SIG_out_norm_7_port, 
      SIG_out_norm_6_port, SIG_out_norm_5_port, SIG_out_norm_4_port, 
      SIG_out_norm_3_port, SIG_out_norm_2_port, EXP_out_norm_7_port, 
      EXP_out_norm_6_port, EXP_out_norm_5_port, EXP_out_norm_4_port, 
      EXP_out_norm_3_port, EXP_out_norm_2_port, EXP_out_norm_1_port, 
      EXP_out_norm_0_port, n91, n92, n93, n94, n_2499, n_2500, n_2501, n_2502, 
      n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510 : 
      std_logic;

begin
   
   SIG_out_norm_27_port <= '0';
   n91 <= '0';
   n92 <= '0';
   n93 <= '0';
   n94 <= '0';
   I9 : FPnormalize_SIG_width28_0 port map( SIG_in(27) => SIG_in(27), 
                           SIG_in(26) => SIG_in(26), SIG_in(25) => SIG_in(25), 
                           SIG_in(24) => SIG_in(24), SIG_in(23) => SIG_in(23), 
                           SIG_in(22) => SIG_in(22), SIG_in(21) => SIG_in(21), 
                           SIG_in(20) => SIG_in(20), SIG_in(19) => SIG_in(19), 
                           SIG_in(18) => SIG_in(18), SIG_in(17) => SIG_in(17), 
                           SIG_in(16) => SIG_in(16), SIG_in(15) => SIG_in(15), 
                           SIG_in(14) => SIG_in(14), SIG_in(13) => SIG_in(13), 
                           SIG_in(12) => SIG_in(12), SIG_in(11) => SIG_in(11), 
                           SIG_in(10) => SIG_in(10), SIG_in(9) => SIG_in(9), 
                           SIG_in(8) => SIG_in(8), SIG_in(7) => SIG_in(7), 
                           SIG_in(6) => SIG_in(6), SIG_in(5) => SIG_in(5), 
                           SIG_in(4) => SIG_in(4), SIG_in(3) => SIG_in(3), 
                           SIG_in(2) => SIG_in(2), SIG_in(1) => n91, SIG_in(0) 
                           => n92, EXP_in(7) => EXP_in(7), EXP_in(6) => 
                           EXP_in(6), EXP_in(5) => EXP_in(5), EXP_in(4) => 
                           EXP_in(4), EXP_in(3) => EXP_in(3), EXP_in(2) => 
                           EXP_in(2), EXP_in(1) => EXP_in(1), EXP_in(0) => 
                           EXP_in(0), SIG_out(27) => n_2499, SIG_out(26) => 
                           SIG_out_norm_26_port, SIG_out(25) => 
                           SIG_out_norm_25_port, SIG_out(24) => 
                           SIG_out_norm_24_port, SIG_out(23) => 
                           SIG_out_norm_23_port, SIG_out(22) => 
                           SIG_out_norm_22_port, SIG_out(21) => 
                           SIG_out_norm_21_port, SIG_out(20) => 
                           SIG_out_norm_20_port, SIG_out(19) => 
                           SIG_out_norm_19_port, SIG_out(18) => 
                           SIG_out_norm_18_port, SIG_out(17) => 
                           SIG_out_norm_17_port, SIG_out(16) => 
                           SIG_out_norm_16_port, SIG_out(15) => 
                           SIG_out_norm_15_port, SIG_out(14) => 
                           SIG_out_norm_14_port, SIG_out(13) => 
                           SIG_out_norm_13_port, SIG_out(12) => 
                           SIG_out_norm_12_port, SIG_out(11) => 
                           SIG_out_norm_11_port, SIG_out(10) => 
                           SIG_out_norm_10_port, SIG_out(9) => 
                           SIG_out_norm_9_port, SIG_out(8) => 
                           SIG_out_norm_8_port, SIG_out(7) => 
                           SIG_out_norm_7_port, SIG_out(6) => 
                           SIG_out_norm_6_port, SIG_out(5) => 
                           SIG_out_norm_5_port, SIG_out(4) => 
                           SIG_out_norm_4_port, SIG_out(3) => 
                           SIG_out_norm_3_port, SIG_out(2) => 
                           SIG_out_norm_2_port, SIG_out(1) => n_2500, 
                           SIG_out(0) => n_2501, EXP_out(7) => 
                           EXP_out_norm_7_port, EXP_out(6) => 
                           EXP_out_norm_6_port, EXP_out(5) => 
                           EXP_out_norm_5_port, EXP_out(4) => 
                           EXP_out_norm_4_port, EXP_out(3) => 
                           EXP_out_norm_3_port, EXP_out(2) => 
                           EXP_out_norm_2_port, EXP_out(1) => 
                           EXP_out_norm_1_port, EXP_out(0) => 
                           EXP_out_norm_0_port, clk => clk);
   I11 : FPround_SIG_width28 port map( SIG_in(27) => SIG_out_norm_27_port, 
                           SIG_in(26) => SIG_out_norm_26_port, SIG_in(25) => 
                           SIG_out_norm_25_port, SIG_in(24) => 
                           SIG_out_norm_24_port, SIG_in(23) => 
                           SIG_out_norm_23_port, SIG_in(22) => 
                           SIG_out_norm_22_port, SIG_in(21) => 
                           SIG_out_norm_21_port, SIG_in(20) => 
                           SIG_out_norm_20_port, SIG_in(19) => 
                           SIG_out_norm_19_port, SIG_in(18) => 
                           SIG_out_norm_18_port, SIG_in(17) => 
                           SIG_out_norm_17_port, SIG_in(16) => 
                           SIG_out_norm_16_port, SIG_in(15) => 
                           SIG_out_norm_15_port, SIG_in(14) => 
                           SIG_out_norm_14_port, SIG_in(13) => 
                           SIG_out_norm_13_port, SIG_in(12) => 
                           SIG_out_norm_12_port, SIG_in(11) => 
                           SIG_out_norm_11_port, SIG_in(10) => 
                           SIG_out_norm_10_port, SIG_in(9) => 
                           SIG_out_norm_9_port, SIG_in(8) => 
                           SIG_out_norm_8_port, SIG_in(7) => 
                           SIG_out_norm_7_port, SIG_in(6) => 
                           SIG_out_norm_6_port, SIG_in(5) => 
                           SIG_out_norm_5_port, SIG_in(4) => 
                           SIG_out_norm_4_port, SIG_in(3) => 
                           SIG_out_norm_3_port, SIG_in(2) => 
                           SIG_out_norm_2_port, SIG_in(1) => n93, SIG_in(0) => 
                           n94, EXP_in(7) => EXP_out_norm_7_port, EXP_in(6) => 
                           EXP_out_norm_6_port, EXP_in(5) => 
                           EXP_out_norm_5_port, EXP_in(4) => 
                           EXP_out_norm_4_port, EXP_in(3) => 
                           EXP_out_norm_3_port, EXP_in(2) => 
                           EXP_out_norm_2_port, EXP_in(1) => 
                           EXP_out_norm_1_port, EXP_in(0) => 
                           EXP_out_norm_0_port, SIG_out(27) => 
                           SIG_out_round(27), SIG_out(26) => SIG_out_round(26),
                           SIG_out(25) => SIG_out_round(25), SIG_out(24) => 
                           SIG_out_round(24), SIG_out(23) => SIG_out_round(23),
                           SIG_out(22) => SIG_out_round(22), SIG_out(21) => 
                           SIG_out_round(21), SIG_out(20) => SIG_out_round(20),
                           SIG_out(19) => SIG_out_round(19), SIG_out(18) => 
                           SIG_out_round(18), SIG_out(17) => SIG_out_round(17),
                           SIG_out(16) => SIG_out_round(16), SIG_out(15) => 
                           SIG_out_round(15), SIG_out(14) => SIG_out_round(14),
                           SIG_out(13) => SIG_out_round(13), SIG_out(12) => 
                           SIG_out_round(12), SIG_out(11) => SIG_out_round(11),
                           SIG_out(10) => SIG_out_round(10), SIG_out(9) => 
                           SIG_out_round(9), SIG_out(8) => SIG_out_round(8), 
                           SIG_out(7) => SIG_out_round(7), SIG_out(6) => 
                           SIG_out_round(6), SIG_out(5) => SIG_out_round(5), 
                           SIG_out(4) => SIG_out_round(4), SIG_out(3) => 
                           SIG_out_round(3), SIG_out(2) => n_2502, SIG_out(1) 
                           => n_2503, SIG_out(0) => n_2504, EXP_out(7) => 
                           EXP_out_round(7), EXP_out(6) => EXP_out_round(6), 
                           EXP_out(5) => EXP_out_round(5), EXP_out(4) => 
                           EXP_out_round(4), EXP_out(3) => EXP_out_round(3), 
                           EXP_out(2) => EXP_out_round(2), EXP_out(1) => 
                           EXP_out_round(1), EXP_out(0) => EXP_out_round(0), 
                           clk => clk);
   MY_CLK_r_REG240_S2 : DFF_X1 port map( D => EXP_pos_stage2, CK => clk, Q => 
                           EXP_pos, QN => n_2505);
   MY_CLK_r_REG237_S2 : DFF_X1 port map( D => EXP_neg_stage2, CK => clk, Q => 
                           EXP_neg, QN => n_2506);
   MY_CLK_r_REG13_S2 : DFF_X1 port map( D => isINF_stage2, CK => clk, Q => 
                           isINF_tab, QN => n_2507);
   MY_CLK_r_REG9_S2 : DFF_X1 port map( D => isZ_tab_stage2, CK => clk, Q => 
                           isZ_tab, QN => n_2508);
   MY_CLK_r_REG5_S2 : DFF_X1 port map( D => isNaN_stage2, CK => clk, Q => isNaN
                           , QN => n_2509);
   MY_CLK_r_REG1_S2 : DFF_X1 port map( D => SIGN_out_stage2, CK => clk, Q => 
                           SIGN_out, QN => n_2510);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage2 is

   port( A_EXP : in std_logic_vector (7 downto 0);  A_SIG : in std_logic_vector
         (31 downto 0);  B_EXP : in std_logic_vector (7 downto 0);  B_SIG : in 
         std_logic_vector (31 downto 0);  SIGN_out_stage1, clk, isINF_stage1, 
         isNaN_stage1, isZ_tab_stage1 : in std_logic;  EXP_in : out 
         std_logic_vector (7 downto 0);  EXP_neg_stage2, EXP_pos_stage2, 
         SIGN_out_stage2 : out std_logic;  SIG_in : out std_logic_vector (27 
         downto 0);  isINF_stage2, isNaN_stage2, isZ_tab_stage2 : out std_logic
         );

end FPmul_stage2;

architecture SYN_struct of FPmul_stage2 is

   component FPmul_stage2_DW01_add_0
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component MBE
      port( A, B : in std_logic_vector (31 downto 0);  C : out std_logic_vector
            (63 downto 0);  clk : in std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic1_port, n130, n131, n132, n133, n134, n135, n136, n137, n139, 
      n140, n141, n142, n143, n144, n145, n146, n120, n121, n122, n123, n124, 
      n125, n126, n127, mw_I4sum_7_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n31, n32, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, 
      n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, 
      n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, 
      n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, 
      n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, 
      n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, 
      n_2581 : std_logic;

begin
   
   X_Logic1_port <= '1';
   U3 : AND2_X1 port map( A1 => n32, A2 => n31, ZN => EXP_pos_stage2);
   U4 : NAND4_X1 port map( A1 => B_EXP(5), A2 => B_EXP(6), A3 => B_EXP(3), A4 
                           => B_EXP(4), ZN => n4);
   U5 : INV_X1 port map( A => B_EXP(0), ZN => n3);
   U6 : INV_X1 port map( A => B_EXP(2), ZN => n2);
   U7 : INV_X1 port map( A => B_EXP(1), ZN => n1);
   U8 : NOR4_X1 port map( A1 => n4, A2 => n3, A3 => n2, A4 => n1, ZN => n10);
   U9 : NAND4_X1 port map( A1 => A_EXP(5), A2 => A_EXP(6), A3 => A_EXP(3), A4 
                           => A_EXP(4), ZN => n8);
   U10 : INV_X1 port map( A => A_EXP(0), ZN => n7);
   U11 : INV_X1 port map( A => A_EXP(2), ZN => n6);
   U12 : INV_X1 port map( A => A_EXP(1), ZN => n5);
   U13 : NOR4_X1 port map( A1 => n8, A2 => n7, A3 => n6, A4 => n5, ZN => n9);
   U14 : NOR4_X1 port map( A1 => B_EXP(7), A2 => A_EXP(7), A3 => n10, A4 => n9,
                           ZN => n127);
   U15 : INV_X1 port map( A => mw_I4sum_7_port, ZN => EXP_in(7));
   MY_CLK_r_REG246_S1 : DFF_X1 port map( D => n120, CK => clk, Q => EXP_in(6), 
                           QN => n_2529);
   MY_CLK_r_REG249_S1 : DFF_X1 port map( D => n121, CK => clk, Q => EXP_in(5), 
                           QN => n_2530);
   MY_CLK_r_REG252_S1 : DFF_X1 port map( D => n122, CK => clk, Q => EXP_in(4), 
                           QN => n_2531);
   MY_CLK_r_REG255_S1 : DFF_X1 port map( D => n123, CK => clk, Q => EXP_in(3), 
                           QN => n_2532);
   MY_CLK_r_REG258_S1 : DFF_X1 port map( D => n124, CK => clk, Q => EXP_in(2), 
                           QN => n_2533);
   MY_CLK_r_REG261_S1 : DFF_X1 port map( D => n125, CK => clk, Q => EXP_in(1), 
                           QN => n_2534);
   MY_CLK_r_REG263_S1 : DFF_X1 port map( D => n126, CK => clk, Q => EXP_in(0), 
                           QN => n_2535);
   MY_CLK_r_REG235_S1 : DFF_X1 port map( D => A_EXP(7), CK => clk, Q => n32, QN
                           => n_2536);
   MY_CLK_r_REG477_S1 : DFF_X1 port map( D => B_EXP(7), CK => clk, Q => n31, QN
                           => n_2537);
   MY_CLK_r_REG0_S1 : DFF_X1 port map( D => SIGN_out_stage1, CK => clk, Q => 
                           SIGN_out_stage2, QN => n_2538);
   MY_CLK_r_REG12_S1 : DFF_X1 port map( D => isINF_stage1, CK => clk, Q => 
                           isINF_stage2, QN => n_2539);
   MY_CLK_r_REG4_S1 : DFF_X1 port map( D => isNaN_stage1, CK => clk, Q => 
                           isNaN_stage2, QN => n_2540);
   MY_CLK_r_REG8_S1 : DFF_X1 port map( D => isZ_tab_stage1, CK => clk, Q => 
                           isZ_tab_stage2, QN => n_2541);
   MY_CLK_r_REG236_S1 : DFF_X1 port map( D => n127, CK => clk, Q => 
                           EXP_neg_stage2, QN => n_2542);
   n146 <= '0';
   n145 <= '0';
   n144 <= '0';
   n143 <= '0';
   n142 <= '0';
   n141 <= '0';
   n140 <= '0';
   n139 <= '0';
   n137 <= '0';
   n136 <= '0';
   n135 <= '0';
   n134 <= '0';
   n133 <= '0';
   n132 <= '0';
   n131 <= '0';
   n130 <= '0';
   MBE_SIG : MBE port map( A(31) => n130, A(30) => n131, A(29) => n132, A(28) 
                           => n133, A(27) => n134, A(26) => n135, A(25) => n136
                           , A(24) => n137, A(23) => A_SIG(23), A(22) => 
                           A_SIG(22), A(21) => A_SIG(21), A(20) => A_SIG(20), 
                           A(19) => A_SIG(19), A(18) => A_SIG(18), A(17) => 
                           A_SIG(17), A(16) => A_SIG(16), A(15) => A_SIG(15), 
                           A(14) => A_SIG(14), A(13) => A_SIG(13), A(12) => 
                           A_SIG(12), A(11) => A_SIG(11), A(10) => A_SIG(10), 
                           A(9) => A_SIG(9), A(8) => A_SIG(8), A(7) => A_SIG(7)
                           , A(6) => A_SIG(6), A(5) => A_SIG(5), A(4) => 
                           A_SIG(4), A(3) => A_SIG(3), A(2) => A_SIG(2), A(1) 
                           => A_SIG(1), A(0) => A_SIG(0), B(31) => n139, B(30) 
                           => n140, B(29) => n141, B(28) => n142, B(27) => n143
                           , B(26) => n144, B(25) => n145, B(24) => n146, B(23)
                           => B_SIG(23), B(22) => B_SIG(22), B(21) => B_SIG(21)
                           , B(20) => B_SIG(20), B(19) => B_SIG(19), B(18) => 
                           B_SIG(18), B(17) => B_SIG(17), B(16) => B_SIG(16), 
                           B(15) => B_SIG(15), B(14) => B_SIG(14), B(13) => 
                           B_SIG(13), B(12) => B_SIG(12), B(11) => B_SIG(11), 
                           B(10) => B_SIG(10), B(9) => B_SIG(9), B(8) => 
                           B_SIG(8), B(7) => B_SIG(7), B(6) => B_SIG(6), B(5) 
                           => B_SIG(5), B(4) => B_SIG(4), B(3) => B_SIG(3), 
                           B(2) => B_SIG(2), B(1) => B_SIG(1), B(0) => B_SIG(0)
                           , C(63) => n_2543, C(62) => n_2544, C(61) => n_2545,
                           C(60) => n_2546, C(59) => n_2547, C(58) => n_2548, 
                           C(57) => n_2549, C(56) => n_2550, C(55) => n_2551, 
                           C(54) => n_2552, C(53) => n_2553, C(52) => n_2554, 
                           C(51) => n_2555, C(50) => n_2556, C(49) => n_2557, 
                           C(48) => n_2558, C(47) => SIG_in(27), C(46) => 
                           SIG_in(26), C(45) => SIG_in(25), C(44) => SIG_in(24)
                           , C(43) => SIG_in(23), C(42) => SIG_in(22), C(41) =>
                           SIG_in(21), C(40) => SIG_in(20), C(39) => SIG_in(19)
                           , C(38) => SIG_in(18), C(37) => SIG_in(17), C(36) =>
                           SIG_in(16), C(35) => SIG_in(15), C(34) => SIG_in(14)
                           , C(33) => SIG_in(13), C(32) => SIG_in(12), C(31) =>
                           SIG_in(11), C(30) => SIG_in(10), C(29) => SIG_in(9),
                           C(28) => SIG_in(8), C(27) => SIG_in(7), C(26) => 
                           SIG_in(6), C(25) => SIG_in(5), C(24) => SIG_in(4), 
                           C(23) => SIG_in(3), C(22) => SIG_in(2), C(21) => 
                           n_2559, C(20) => n_2560, C(19) => n_2561, C(18) => 
                           n_2562, C(17) => n_2563, C(16) => n_2564, C(15) => 
                           n_2565, C(14) => n_2566, C(13) => n_2567, C(12) => 
                           n_2568, C(11) => n_2569, C(10) => n_2570, C(9) => 
                           n_2571, C(8) => n_2572, C(7) => n_2573, C(6) => 
                           n_2574, C(5) => n_2575, C(4) => n_2576, C(3) => 
                           n_2577, C(2) => n_2578, C(1) => n_2579, C(0) => 
                           n_2580, clk => clk);
   add_1_root_add_131_2 : FPmul_stage2_DW01_add_0 port map( A(7) => n32, A(6) 
                           => A_EXP(6), A(5) => A_EXP(5), A(4) => A_EXP(4), 
                           A(3) => A_EXP(3), A(2) => A_EXP(2), A(1) => A_EXP(1)
                           , A(0) => A_EXP(0), B(7) => n31, B(6) => B_EXP(6), 
                           B(5) => B_EXP(5), B(4) => B_EXP(4), B(3) => B_EXP(3)
                           , B(2) => B_EXP(2), B(1) => B_EXP(1), B(0) => 
                           B_EXP(0), CI => X_Logic1_port, SUM(7) => 
                           mw_I4sum_7_port, SUM(6) => n120, SUM(5) => n121, 
                           SUM(4) => n122, SUM(3) => n123, SUM(2) => n124, 
                           SUM(1) => n125, SUM(0) => n126, CO => n_2581, clk =>
                           clk);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage1 is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         A_EXP : out std_logic_vector (7 downto 0);  A_SIG : out 
         std_logic_vector (31 downto 0);  B_EXP : out std_logic_vector (7 
         downto 0);  B_SIG : out std_logic_vector (31 downto 0);  
         SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : out 
         std_logic);

end FPmul_stage1;

architecture SYN_struct of FPmul_stage1 is

   component UnpackFP_1
      port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector
            (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, 
            isNaN, isINF, isZ, isDN : out std_logic);
   end component;
   
   component UnpackFP_0
      port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector
            (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, 
            isNaN, isINF, isZ, isDN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal A_isINF, A_isNaN, A_isZ, B_isINF, B_isNaN, B_isZ, A_SIGN, B_SIGN, n18
      , n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n_2598, n_2599, 
      n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, 
      n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615 : std_logic;

begin
   
   U26 : INV_X1 port map( A => B_isZ, ZN => n20);
   U27 : INV_X1 port map( A => A_isZ, ZN => n22);
   U28 : OR2_X1 port map( A1 => B_isNaN, A2 => A_isNaN, ZN => n21);
   U29 : INV_X1 port map( A => n21, ZN => n18);
   U30 : INV_X1 port map( A => A_isINF, ZN => n25);
   U31 : NAND2_X1 port map( A1 => n18, A2 => n25, ZN => n19);
   U32 : AOI211_X1 port map( C1 => n20, C2 => n22, A => n19, B => B_isINF, ZN 
                           => isZ_tab_stage1);
   U33 : NAND2_X1 port map( A1 => B_isZ, A2 => A_isINF, ZN => n26);
   U34 : NAND2_X1 port map( A1 => n21, A2 => n25, ZN => n23);
   U35 : MUX2_X1 port map( A => n23, B => n22, S => B_isINF, Z => n24);
   U36 : NAND2_X1 port map( A1 => n26, A2 => n24, ZN => isNaN_stage1);
   U37 : NOR2_X1 port map( A1 => B_isZ, A2 => n25, ZN => n29);
   U38 : INV_X1 port map( A => n26, ZN => n27);
   U39 : NOR2_X1 port map( A1 => A_isZ, A2 => n27, ZN => n28);
   U40 : MUX2_X1 port map( A => n29, B => n28, S => B_isINF, Z => isINF_stage1)
                           ;
   U41 : XOR2_X1 port map( A => B_SIGN, B => A_SIGN, Z => SIGN_out_stage1);
   I0 : UnpackFP_0 port map( FP(31) => FP_A(31), FP(30) => FP_A(30), FP(29) => 
                           FP_A(29), FP(28) => FP_A(28), FP(27) => FP_A(27), 
                           FP(26) => FP_A(26), FP(25) => FP_A(25), FP(24) => 
                           FP_A(24), FP(23) => FP_A(23), FP(22) => FP_A(22), 
                           FP(21) => FP_A(21), FP(20) => FP_A(20), FP(19) => 
                           FP_A(19), FP(18) => FP_A(18), FP(17) => FP_A(17), 
                           FP(16) => FP_A(16), FP(15) => FP_A(15), FP(14) => 
                           FP_A(14), FP(13) => FP_A(13), FP(12) => FP_A(12), 
                           FP(11) => FP_A(11), FP(10) => FP_A(10), FP(9) => 
                           FP_A(9), FP(8) => FP_A(8), FP(7) => FP_A(7), FP(6) 
                           => FP_A(6), FP(5) => FP_A(5), FP(4) => FP_A(4), 
                           FP(3) => FP_A(3), FP(2) => FP_A(2), FP(1) => FP_A(1)
                           , FP(0) => FP_A(0), SIG(31) => n_2598, SIG(30) => 
                           n_2599, SIG(29) => n_2600, SIG(28) => n_2601, 
                           SIG(27) => n_2602, SIG(26) => n_2603, SIG(25) => 
                           n_2604, SIG(24) => n_2605, SIG(23) => A_SIG(23), 
                           SIG(22) => A_SIG(22), SIG(21) => A_SIG(21), SIG(20) 
                           => A_SIG(20), SIG(19) => A_SIG(19), SIG(18) => 
                           A_SIG(18), SIG(17) => A_SIG(17), SIG(16) => 
                           A_SIG(16), SIG(15) => A_SIG(15), SIG(14) => 
                           A_SIG(14), SIG(13) => A_SIG(13), SIG(12) => 
                           A_SIG(12), SIG(11) => A_SIG(11), SIG(10) => 
                           A_SIG(10), SIG(9) => A_SIG(9), SIG(8) => A_SIG(8), 
                           SIG(7) => A_SIG(7), SIG(6) => A_SIG(6), SIG(5) => 
                           A_SIG(5), SIG(4) => A_SIG(4), SIG(3) => A_SIG(3), 
                           SIG(2) => A_SIG(2), SIG(1) => A_SIG(1), SIG(0) => 
                           A_SIG(0), EXP(7) => A_EXP(7), EXP(6) => A_EXP(6), 
                           EXP(5) => A_EXP(5), EXP(4) => A_EXP(4), EXP(3) => 
                           A_EXP(3), EXP(2) => A_EXP(2), EXP(1) => A_EXP(1), 
                           EXP(0) => A_EXP(0), SIGN => A_SIGN, isNaN => A_isNaN
                           , isINF => A_isINF, isZ => A_isZ, isDN => n_2606);
   I1 : UnpackFP_1 port map( FP(31) => FP_B(31), FP(30) => FP_B(30), FP(29) => 
                           FP_B(29), FP(28) => FP_B(28), FP(27) => FP_B(27), 
                           FP(26) => FP_B(26), FP(25) => FP_B(25), FP(24) => 
                           FP_B(24), FP(23) => FP_B(23), FP(22) => FP_B(22), 
                           FP(21) => FP_B(21), FP(20) => FP_B(20), FP(19) => 
                           FP_B(19), FP(18) => FP_B(18), FP(17) => FP_B(17), 
                           FP(16) => FP_B(16), FP(15) => FP_B(15), FP(14) => 
                           FP_B(14), FP(13) => FP_B(13), FP(12) => FP_B(12), 
                           FP(11) => FP_B(11), FP(10) => FP_B(10), FP(9) => 
                           FP_B(9), FP(8) => FP_B(8), FP(7) => FP_B(7), FP(6) 
                           => FP_B(6), FP(5) => FP_B(5), FP(4) => FP_B(4), 
                           FP(3) => FP_B(3), FP(2) => FP_B(2), FP(1) => FP_B(1)
                           , FP(0) => FP_B(0), SIG(31) => n_2607, SIG(30) => 
                           n_2608, SIG(29) => n_2609, SIG(28) => n_2610, 
                           SIG(27) => n_2611, SIG(26) => n_2612, SIG(25) => 
                           n_2613, SIG(24) => n_2614, SIG(23) => B_SIG(23), 
                           SIG(22) => B_SIG(22), SIG(21) => B_SIG(21), SIG(20) 
                           => B_SIG(20), SIG(19) => B_SIG(19), SIG(18) => 
                           B_SIG(18), SIG(17) => B_SIG(17), SIG(16) => 
                           B_SIG(16), SIG(15) => B_SIG(15), SIG(14) => 
                           B_SIG(14), SIG(13) => B_SIG(13), SIG(12) => 
                           B_SIG(12), SIG(11) => B_SIG(11), SIG(10) => 
                           B_SIG(10), SIG(9) => B_SIG(9), SIG(8) => B_SIG(8), 
                           SIG(7) => B_SIG(7), SIG(6) => B_SIG(6), SIG(5) => 
                           B_SIG(5), SIG(4) => B_SIG(4), SIG(3) => B_SIG(3), 
                           SIG(2) => B_SIG(2), SIG(1) => B_SIG(1), SIG(0) => 
                           B_SIG(0), EXP(7) => B_EXP(7), EXP(6) => B_EXP(6), 
                           EXP(5) => B_EXP(5), EXP(4) => B_EXP(4), EXP(3) => 
                           B_EXP(3), EXP(2) => B_EXP(2), EXP(1) => B_EXP(1), 
                           EXP(0) => B_EXP(0), SIGN => B_SIGN, isNaN => B_isNaN
                           , isINF => B_isINF, isZ => B_isZ, isDN => n_2615);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         FP_Z : out std_logic_vector (31 downto 0));

end FPmul;

architecture SYN_pipeline of FPmul is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FPmul_stage4
      port( EXP_neg : in std_logic;  EXP_out_round : in std_logic_vector (7 
            downto 0);  EXP_pos, SIGN_out : in std_logic;  SIG_out_round : in 
            std_logic_vector (27 downto 0);  clk, isINF_tab, isNaN, isZ_tab : 
            in std_logic;  FP_Z : out std_logic_vector (31 downto 0));
   end component;
   
   component FPmul_stage3
      port( EXP_in : in std_logic_vector (7 downto 0);  EXP_neg_stage2, 
            EXP_pos_stage2, SIGN_out_stage2 : in std_logic;  SIG_in : in 
            std_logic_vector (27 downto 0);  clk, isINF_stage2, isNaN_stage2, 
            isZ_tab_stage2 : in std_logic;  EXP_neg : out std_logic;  
            EXP_out_round : out std_logic_vector (7 downto 0);  EXP_pos, 
            SIGN_out : out std_logic;  SIG_out_round : out std_logic_vector (27
            downto 0);  isINF_tab, isNaN, isZ_tab : out std_logic);
   end component;
   
   component FPmul_stage2
      port( A_EXP : in std_logic_vector (7 downto 0);  A_SIG : in 
            std_logic_vector (31 downto 0);  B_EXP : in std_logic_vector (7 
            downto 0);  B_SIG : in std_logic_vector (31 downto 0);  
            SIGN_out_stage1, clk, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : 
            in std_logic;  EXP_in : out std_logic_vector (7 downto 0);  
            EXP_neg_stage2, EXP_pos_stage2, SIGN_out_stage2 : out std_logic;  
            SIG_in : out std_logic_vector (27 downto 0);  isINF_stage2, 
            isNaN_stage2, isZ_tab_stage2 : out std_logic);
   end component;
   
   component FPmul_stage1
      port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic
            ;  A_EXP : out std_logic_vector (7 downto 0);  A_SIG : out 
            std_logic_vector (31 downto 0);  B_EXP : out std_logic_vector (7 
            downto 0);  B_SIG : out std_logic_vector (31 downto 0);  
            SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : out 
            std_logic);
   end component;
   
   signal n8, A_EXP_7_port, A_EXP_6_port, A_EXP_5_port, A_EXP_4_port, 
      A_EXP_3_port, A_EXP_2_port, A_EXP_1_port, A_EXP_0_port, A_SIG_22_port, 
      A_SIG_21_port, A_SIG_20_port, A_SIG_19_port, A_SIG_18_port, A_SIG_17_port
      , A_SIG_16_port, A_SIG_15_port, A_SIG_14_port, A_SIG_13_port, 
      A_SIG_12_port, A_SIG_11_port, A_SIG_10_port, A_SIG_9_port, A_SIG_8_port, 
      A_SIG_7_port, A_SIG_6_port, A_SIG_5_port, A_SIG_4_port, A_SIG_3_port, 
      A_SIG_2_port, A_SIG_1_port, A_SIG_0_port, B_EXP_7_port, B_EXP_6_port, 
      B_EXP_5_port, B_EXP_4_port, B_EXP_3_port, B_EXP_2_port, B_EXP_1_port, 
      B_EXP_0_port, B_SIG_22_port, B_SIG_21_port, B_SIG_20_port, B_SIG_19_port,
      B_SIG_18_port, B_SIG_17_port, B_SIG_16_port, B_SIG_15_port, B_SIG_14_port
      , B_SIG_13_port, B_SIG_12_port, B_SIG_11_port, B_SIG_10_port, 
      B_SIG_9_port, B_SIG_8_port, B_SIG_7_port, B_SIG_6_port, B_SIG_5_port, 
      B_SIG_4_port, B_SIG_3_port, B_SIG_2_port, B_SIG_1_port, B_SIG_0_port, 
      SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1, 
      EXP_in_7_port, EXP_in_6_port, EXP_in_5_port, EXP_in_4_port, EXP_in_3_port
      , EXP_in_2_port, EXP_in_1_port, EXP_in_0_port, EXP_neg_stage2, 
      EXP_pos_stage2, SIGN_out_stage2, SIG_in_27_port, SIG_in_26_port, 
      SIG_in_25_port, SIG_in_24_port, SIG_in_23_port, SIG_in_22_port, 
      SIG_in_21_port, SIG_in_20_port, SIG_in_19_port, SIG_in_18_port, 
      SIG_in_17_port, SIG_in_16_port, SIG_in_15_port, SIG_in_14_port, 
      SIG_in_13_port, SIG_in_12_port, SIG_in_11_port, SIG_in_10_port, 
      SIG_in_9_port, SIG_in_8_port, SIG_in_7_port, SIG_in_6_port, SIG_in_5_port
      , SIG_in_4_port, SIG_in_3_port, SIG_in_2_port, isINF_stage2, isNaN_stage2
      , isZ_tab_stage2, EXP_neg, EXP_out_round_7_port, EXP_out_round_6_port, 
      EXP_out_round_5_port, EXP_out_round_4_port, EXP_out_round_3_port, 
      EXP_out_round_2_port, EXP_out_round_1_port, EXP_out_round_0_port, EXP_pos
      , SIGN_out, SIG_out_round_26_port, SIG_out_round_25_port, 
      SIG_out_round_24_port, SIG_out_round_23_port, SIG_out_round_22_port, 
      SIG_out_round_21_port, SIG_out_round_20_port, SIG_out_round_19_port, 
      SIG_out_round_18_port, SIG_out_round_17_port, SIG_out_round_16_port, 
      SIG_out_round_15_port, SIG_out_round_14_port, SIG_out_round_13_port, 
      SIG_out_round_12_port, SIG_out_round_11_port, SIG_out_round_10_port, 
      SIG_out_round_9_port, SIG_out_round_8_port, SIG_out_round_7_port, 
      SIG_out_round_6_port, SIG_out_round_5_port, SIG_out_round_4_port, 
      SIG_out_round_3_port, isINF_tab, isNaN, isZ_tab, n1, n4, n5, n6, n7, n9, 
      n10, n12, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623,
      n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, 
      n_2633, n_2634, n_2635, n_2636, n_2637 : std_logic;

begin
   
   n1 <= '0';
   n4 <= '0';
   n5 <= '0';
   n6 <= '0';
   n7 <= '0';
   I1 : FPmul_stage1 port map( FP_A(31) => FP_A(31), FP_A(30) => FP_A(30), 
                           FP_A(29) => FP_A(29), FP_A(28) => FP_A(28), FP_A(27)
                           => FP_A(27), FP_A(26) => FP_A(26), FP_A(25) => 
                           FP_A(25), FP_A(24) => FP_A(24), FP_A(23) => FP_A(23)
                           , FP_A(22) => FP_A(22), FP_A(21) => FP_A(21), 
                           FP_A(20) => FP_A(20), FP_A(19) => FP_A(19), FP_A(18)
                           => FP_A(18), FP_A(17) => FP_A(17), FP_A(16) => 
                           FP_A(16), FP_A(15) => FP_A(15), FP_A(14) => FP_A(14)
                           , FP_A(13) => FP_A(13), FP_A(12) => FP_A(12), 
                           FP_A(11) => FP_A(11), FP_A(10) => FP_A(10), FP_A(9) 
                           => FP_A(9), FP_A(8) => FP_A(8), FP_A(7) => FP_A(7), 
                           FP_A(6) => FP_A(6), FP_A(5) => FP_A(5), FP_A(4) => 
                           FP_A(4), FP_A(3) => FP_A(3), FP_A(2) => FP_A(2), 
                           FP_A(1) => FP_A(1), FP_A(0) => FP_A(0), FP_B(31) => 
                           FP_B(31), FP_B(30) => FP_B(30), FP_B(29) => FP_B(29)
                           , FP_B(28) => FP_B(28), FP_B(27) => FP_B(27), 
                           FP_B(26) => FP_B(26), FP_B(25) => FP_B(25), FP_B(24)
                           => FP_B(24), FP_B(23) => FP_B(23), FP_B(22) => 
                           FP_B(22), FP_B(21) => FP_B(21), FP_B(20) => FP_B(20)
                           , FP_B(19) => FP_B(19), FP_B(18) => FP_B(18), 
                           FP_B(17) => FP_B(17), FP_B(16) => FP_B(16), FP_B(15)
                           => FP_B(15), FP_B(14) => FP_B(14), FP_B(13) => 
                           FP_B(13), FP_B(12) => FP_B(12), FP_B(11) => FP_B(11)
                           , FP_B(10) => FP_B(10), FP_B(9) => FP_B(9), FP_B(8) 
                           => FP_B(8), FP_B(7) => FP_B(7), FP_B(6) => FP_B(6), 
                           FP_B(5) => FP_B(5), FP_B(4) => FP_B(4), FP_B(3) => 
                           FP_B(3), FP_B(2) => FP_B(2), FP_B(1) => FP_B(1), 
                           FP_B(0) => FP_B(0), clk => clk, A_EXP(7) => 
                           A_EXP_7_port, A_EXP(6) => A_EXP_6_port, A_EXP(5) => 
                           A_EXP_5_port, A_EXP(4) => A_EXP_4_port, A_EXP(3) => 
                           A_EXP_3_port, A_EXP(2) => A_EXP_2_port, A_EXP(1) => 
                           A_EXP_1_port, A_EXP(0) => A_EXP_0_port, A_SIG(31) =>
                           n_2616, A_SIG(30) => n_2617, A_SIG(29) => n_2618, 
                           A_SIG(28) => n_2619, A_SIG(27) => n_2620, A_SIG(26) 
                           => n_2621, A_SIG(25) => n_2622, A_SIG(24) => n_2623,
                           A_SIG(23) => n12, A_SIG(22) => A_SIG_22_port, 
                           A_SIG(21) => A_SIG_21_port, A_SIG(20) => 
                           A_SIG_20_port, A_SIG(19) => A_SIG_19_port, A_SIG(18)
                           => A_SIG_18_port, A_SIG(17) => A_SIG_17_port, 
                           A_SIG(16) => A_SIG_16_port, A_SIG(15) => 
                           A_SIG_15_port, A_SIG(14) => A_SIG_14_port, A_SIG(13)
                           => A_SIG_13_port, A_SIG(12) => A_SIG_12_port, 
                           A_SIG(11) => A_SIG_11_port, A_SIG(10) => 
                           A_SIG_10_port, A_SIG(9) => A_SIG_9_port, A_SIG(8) =>
                           A_SIG_8_port, A_SIG(7) => A_SIG_7_port, A_SIG(6) => 
                           A_SIG_6_port, A_SIG(5) => A_SIG_5_port, A_SIG(4) => 
                           A_SIG_4_port, A_SIG(3) => A_SIG_3_port, A_SIG(2) => 
                           A_SIG_2_port, A_SIG(1) => A_SIG_1_port, A_SIG(0) => 
                           A_SIG_0_port, B_EXP(7) => B_EXP_7_port, B_EXP(6) => 
                           B_EXP_6_port, B_EXP(5) => B_EXP_5_port, B_EXP(4) => 
                           B_EXP_4_port, B_EXP(3) => B_EXP_3_port, B_EXP(2) => 
                           B_EXP_2_port, B_EXP(1) => B_EXP_1_port, B_EXP(0) => 
                           B_EXP_0_port, B_SIG(31) => n_2624, B_SIG(30) => 
                           n_2625, B_SIG(29) => n_2626, B_SIG(28) => n_2627, 
                           B_SIG(27) => n_2628, B_SIG(26) => n_2629, B_SIG(25) 
                           => n_2630, B_SIG(24) => n_2631, B_SIG(23) => n10, 
                           B_SIG(22) => B_SIG_22_port, B_SIG(21) => 
                           B_SIG_21_port, B_SIG(20) => B_SIG_20_port, B_SIG(19)
                           => B_SIG_19_port, B_SIG(18) => B_SIG_18_port, 
                           B_SIG(17) => B_SIG_17_port, B_SIG(16) => 
                           B_SIG_16_port, B_SIG(15) => B_SIG_15_port, B_SIG(14)
                           => B_SIG_14_port, B_SIG(13) => B_SIG_13_port, 
                           B_SIG(12) => B_SIG_12_port, B_SIG(11) => 
                           B_SIG_11_port, B_SIG(10) => B_SIG_10_port, B_SIG(9) 
                           => B_SIG_9_port, B_SIG(8) => B_SIG_8_port, B_SIG(7) 
                           => B_SIG_7_port, B_SIG(6) => B_SIG_6_port, B_SIG(5) 
                           => B_SIG_5_port, B_SIG(4) => B_SIG_4_port, B_SIG(3) 
                           => B_SIG_3_port, B_SIG(2) => B_SIG_2_port, B_SIG(1) 
                           => B_SIG_1_port, B_SIG(0) => B_SIG_0_port, 
                           SIGN_out_stage1 => SIGN_out_stage1, isINF_stage1 => 
                           isINF_stage1, isNaN_stage1 => isNaN_stage1, 
                           isZ_tab_stage1 => isZ_tab_stage1);
   I2 : FPmul_stage2 port map( A_EXP(7) => A_EXP_7_port, A_EXP(6) => 
                           A_EXP_6_port, A_EXP(5) => A_EXP_5_port, A_EXP(4) => 
                           A_EXP_4_port, A_EXP(3) => A_EXP_3_port, A_EXP(2) => 
                           A_EXP_2_port, A_EXP(1) => A_EXP_1_port, A_EXP(0) => 
                           A_EXP_0_port, A_SIG(31) => n1, A_SIG(30) => n1, 
                           A_SIG(29) => n1, A_SIG(28) => n1, A_SIG(27) => n1, 
                           A_SIG(26) => n1, A_SIG(25) => n1, A_SIG(24) => n1, 
                           A_SIG(23) => n12, A_SIG(22) => A_SIG_22_port, 
                           A_SIG(21) => A_SIG_21_port, A_SIG(20) => 
                           A_SIG_20_port, A_SIG(19) => A_SIG_19_port, A_SIG(18)
                           => A_SIG_18_port, A_SIG(17) => A_SIG_17_port, 
                           A_SIG(16) => A_SIG_16_port, A_SIG(15) => 
                           A_SIG_15_port, A_SIG(14) => A_SIG_14_port, A_SIG(13)
                           => A_SIG_13_port, A_SIG(12) => A_SIG_12_port, 
                           A_SIG(11) => A_SIG_11_port, A_SIG(10) => 
                           A_SIG_10_port, A_SIG(9) => A_SIG_9_port, A_SIG(8) =>
                           A_SIG_8_port, A_SIG(7) => A_SIG_7_port, A_SIG(6) => 
                           A_SIG_6_port, A_SIG(5) => A_SIG_5_port, A_SIG(4) => 
                           A_SIG_4_port, A_SIG(3) => A_SIG_3_port, A_SIG(2) => 
                           A_SIG_2_port, A_SIG(1) => A_SIG_1_port, A_SIG(0) => 
                           A_SIG_0_port, B_EXP(7) => B_EXP_7_port, B_EXP(6) => 
                           B_EXP_6_port, B_EXP(5) => B_EXP_5_port, B_EXP(4) => 
                           B_EXP_4_port, B_EXP(3) => B_EXP_3_port, B_EXP(2) => 
                           B_EXP_2_port, B_EXP(1) => B_EXP_1_port, B_EXP(0) => 
                           B_EXP_0_port, B_SIG(31) => n1, B_SIG(30) => n1, 
                           B_SIG(29) => n1, B_SIG(28) => n1, B_SIG(27) => n1, 
                           B_SIG(26) => n1, B_SIG(25) => n1, B_SIG(24) => n1, 
                           B_SIG(23) => n10, B_SIG(22) => B_SIG_22_port, 
                           B_SIG(21) => B_SIG_21_port, B_SIG(20) => 
                           B_SIG_20_port, B_SIG(19) => B_SIG_19_port, B_SIG(18)
                           => B_SIG_18_port, B_SIG(17) => B_SIG_17_port, 
                           B_SIG(16) => B_SIG_16_port, B_SIG(15) => 
                           B_SIG_15_port, B_SIG(14) => B_SIG_14_port, B_SIG(13)
                           => B_SIG_13_port, B_SIG(12) => B_SIG_12_port, 
                           B_SIG(11) => B_SIG_11_port, B_SIG(10) => 
                           B_SIG_10_port, B_SIG(9) => B_SIG_9_port, B_SIG(8) =>
                           B_SIG_8_port, B_SIG(7) => B_SIG_7_port, B_SIG(6) => 
                           B_SIG_6_port, B_SIG(5) => B_SIG_5_port, B_SIG(4) => 
                           B_SIG_4_port, B_SIG(3) => B_SIG_3_port, B_SIG(2) => 
                           B_SIG_2_port, B_SIG(1) => B_SIG_1_port, B_SIG(0) => 
                           B_SIG_0_port, SIGN_out_stage1 => SIGN_out_stage1, 
                           clk => clk, isINF_stage1 => isINF_stage1, 
                           isNaN_stage1 => isNaN_stage1, isZ_tab_stage1 => 
                           isZ_tab_stage1, EXP_in(7) => EXP_in_7_port, 
                           EXP_in(6) => EXP_in_6_port, EXP_in(5) => 
                           EXP_in_5_port, EXP_in(4) => EXP_in_4_port, EXP_in(3)
                           => EXP_in_3_port, EXP_in(2) => EXP_in_2_port, 
                           EXP_in(1) => EXP_in_1_port, EXP_in(0) => 
                           EXP_in_0_port, EXP_neg_stage2 => EXP_neg_stage2, 
                           EXP_pos_stage2 => EXP_pos_stage2, SIGN_out_stage2 =>
                           SIGN_out_stage2, SIG_in(27) => SIG_in_27_port, 
                           SIG_in(26) => SIG_in_26_port, SIG_in(25) => 
                           SIG_in_25_port, SIG_in(24) => SIG_in_24_port, 
                           SIG_in(23) => SIG_in_23_port, SIG_in(22) => 
                           SIG_in_22_port, SIG_in(21) => SIG_in_21_port, 
                           SIG_in(20) => SIG_in_20_port, SIG_in(19) => 
                           SIG_in_19_port, SIG_in(18) => SIG_in_18_port, 
                           SIG_in(17) => SIG_in_17_port, SIG_in(16) => 
                           SIG_in_16_port, SIG_in(15) => SIG_in_15_port, 
                           SIG_in(14) => SIG_in_14_port, SIG_in(13) => 
                           SIG_in_13_port, SIG_in(12) => SIG_in_12_port, 
                           SIG_in(11) => SIG_in_11_port, SIG_in(10) => 
                           SIG_in_10_port, SIG_in(9) => SIG_in_9_port, 
                           SIG_in(8) => SIG_in_8_port, SIG_in(7) => 
                           SIG_in_7_port, SIG_in(6) => SIG_in_6_port, SIG_in(5)
                           => SIG_in_5_port, SIG_in(4) => SIG_in_4_port, 
                           SIG_in(3) => SIG_in_3_port, SIG_in(2) => 
                           SIG_in_2_port, SIG_in(1) => n_2632, SIG_in(0) => 
                           n_2633, isINF_stage2 => isINF_stage2, isNaN_stage2 
                           => isNaN_stage2, isZ_tab_stage2 => isZ_tab_stage2);
   I3 : FPmul_stage3 port map( EXP_in(7) => EXP_in_7_port, EXP_in(6) => 
                           EXP_in_6_port, EXP_in(5) => EXP_in_5_port, EXP_in(4)
                           => EXP_in_4_port, EXP_in(3) => EXP_in_3_port, 
                           EXP_in(2) => EXP_in_2_port, EXP_in(1) => 
                           EXP_in_1_port, EXP_in(0) => EXP_in_0_port, 
                           EXP_neg_stage2 => EXP_neg_stage2, EXP_pos_stage2 => 
                           EXP_pos_stage2, SIGN_out_stage2 => SIGN_out_stage2, 
                           SIG_in(27) => SIG_in_27_port, SIG_in(26) => 
                           SIG_in_26_port, SIG_in(25) => SIG_in_25_port, 
                           SIG_in(24) => SIG_in_24_port, SIG_in(23) => 
                           SIG_in_23_port, SIG_in(22) => SIG_in_22_port, 
                           SIG_in(21) => SIG_in_21_port, SIG_in(20) => 
                           SIG_in_20_port, SIG_in(19) => SIG_in_19_port, 
                           SIG_in(18) => SIG_in_18_port, SIG_in(17) => 
                           SIG_in_17_port, SIG_in(16) => SIG_in_16_port, 
                           SIG_in(15) => SIG_in_15_port, SIG_in(14) => 
                           SIG_in_14_port, SIG_in(13) => SIG_in_13_port, 
                           SIG_in(12) => SIG_in_12_port, SIG_in(11) => 
                           SIG_in_11_port, SIG_in(10) => SIG_in_10_port, 
                           SIG_in(9) => SIG_in_9_port, SIG_in(8) => 
                           SIG_in_8_port, SIG_in(7) => SIG_in_7_port, SIG_in(6)
                           => SIG_in_6_port, SIG_in(5) => SIG_in_5_port, 
                           SIG_in(4) => SIG_in_4_port, SIG_in(3) => 
                           SIG_in_3_port, SIG_in(2) => SIG_in_2_port, SIG_in(1)
                           => n4, SIG_in(0) => n5, clk => clk, isINF_stage2 => 
                           isINF_stage2, isNaN_stage2 => isNaN_stage2, 
                           isZ_tab_stage2 => isZ_tab_stage2, EXP_neg => EXP_neg
                           , EXP_out_round(7) => EXP_out_round_7_port, 
                           EXP_out_round(6) => EXP_out_round_6_port, 
                           EXP_out_round(5) => EXP_out_round_5_port, 
                           EXP_out_round(4) => EXP_out_round_4_port, 
                           EXP_out_round(3) => EXP_out_round_3_port, 
                           EXP_out_round(2) => EXP_out_round_2_port, 
                           EXP_out_round(1) => EXP_out_round_1_port, 
                           EXP_out_round(0) => EXP_out_round_0_port, EXP_pos =>
                           EXP_pos, SIGN_out => SIGN_out, SIG_out_round(27) => 
                           n9, SIG_out_round(26) => SIG_out_round_26_port, 
                           SIG_out_round(25) => SIG_out_round_25_port, 
                           SIG_out_round(24) => SIG_out_round_24_port, 
                           SIG_out_round(23) => SIG_out_round_23_port, 
                           SIG_out_round(22) => SIG_out_round_22_port, 
                           SIG_out_round(21) => SIG_out_round_21_port, 
                           SIG_out_round(20) => SIG_out_round_20_port, 
                           SIG_out_round(19) => SIG_out_round_19_port, 
                           SIG_out_round(18) => SIG_out_round_18_port, 
                           SIG_out_round(17) => SIG_out_round_17_port, 
                           SIG_out_round(16) => SIG_out_round_16_port, 
                           SIG_out_round(15) => SIG_out_round_15_port, 
                           SIG_out_round(14) => SIG_out_round_14_port, 
                           SIG_out_round(13) => SIG_out_round_13_port, 
                           SIG_out_round(12) => SIG_out_round_12_port, 
                           SIG_out_round(11) => SIG_out_round_11_port, 
                           SIG_out_round(10) => SIG_out_round_10_port, 
                           SIG_out_round(9) => SIG_out_round_9_port, 
                           SIG_out_round(8) => SIG_out_round_8_port, 
                           SIG_out_round(7) => SIG_out_round_7_port, 
                           SIG_out_round(6) => SIG_out_round_6_port, 
                           SIG_out_round(5) => SIG_out_round_5_port, 
                           SIG_out_round(4) => SIG_out_round_4_port, 
                           SIG_out_round(3) => SIG_out_round_3_port, 
                           SIG_out_round(2) => n_2634, SIG_out_round(1) => 
                           n_2635, SIG_out_round(0) => n_2636, isINF_tab => 
                           isINF_tab, isNaN => isNaN, isZ_tab => isZ_tab);
   I4 : FPmul_stage4 port map( EXP_neg => EXP_neg, EXP_out_round(7) => 
                           EXP_out_round_7_port, EXP_out_round(6) => 
                           EXP_out_round_6_port, EXP_out_round(5) => 
                           EXP_out_round_5_port, EXP_out_round(4) => 
                           EXP_out_round_4_port, EXP_out_round(3) => 
                           EXP_out_round_3_port, EXP_out_round(2) => 
                           EXP_out_round_2_port, EXP_out_round(1) => 
                           EXP_out_round_1_port, EXP_out_round(0) => 
                           EXP_out_round_0_port, EXP_pos => EXP_pos, SIGN_out 
                           => SIGN_out, SIG_out_round(27) => n9, 
                           SIG_out_round(26) => SIG_out_round_26_port, 
                           SIG_out_round(25) => SIG_out_round_25_port, 
                           SIG_out_round(24) => SIG_out_round_24_port, 
                           SIG_out_round(23) => SIG_out_round_23_port, 
                           SIG_out_round(22) => SIG_out_round_22_port, 
                           SIG_out_round(21) => SIG_out_round_21_port, 
                           SIG_out_round(20) => SIG_out_round_20_port, 
                           SIG_out_round(19) => SIG_out_round_19_port, 
                           SIG_out_round(18) => SIG_out_round_18_port, 
                           SIG_out_round(17) => SIG_out_round_17_port, 
                           SIG_out_round(16) => SIG_out_round_16_port, 
                           SIG_out_round(15) => SIG_out_round_15_port, 
                           SIG_out_round(14) => SIG_out_round_14_port, 
                           SIG_out_round(13) => SIG_out_round_13_port, 
                           SIG_out_round(12) => SIG_out_round_12_port, 
                           SIG_out_round(11) => SIG_out_round_11_port, 
                           SIG_out_round(10) => SIG_out_round_10_port, 
                           SIG_out_round(9) => SIG_out_round_9_port, 
                           SIG_out_round(8) => SIG_out_round_8_port, 
                           SIG_out_round(7) => SIG_out_round_7_port, 
                           SIG_out_round(6) => SIG_out_round_6_port, 
                           SIG_out_round(5) => SIG_out_round_5_port, 
                           SIG_out_round(4) => SIG_out_round_4_port, 
                           SIG_out_round(3) => SIG_out_round_3_port, 
                           SIG_out_round(2) => n1, SIG_out_round(1) => n6, 
                           SIG_out_round(0) => n7, clk => clk, isINF_tab => 
                           isINF_tab, isNaN => isNaN, isZ_tab => isZ_tab, 
                           FP_Z(31) => n8, FP_Z(30) => FP_Z(30), FP_Z(29) => 
                           FP_Z(29), FP_Z(28) => FP_Z(28), FP_Z(27) => FP_Z(27)
                           , FP_Z(26) => FP_Z(26), FP_Z(25) => FP_Z(25), 
                           FP_Z(24) => FP_Z(24), FP_Z(23) => FP_Z(23), FP_Z(22)
                           => FP_Z(22), FP_Z(21) => FP_Z(21), FP_Z(20) => 
                           FP_Z(20), FP_Z(19) => FP_Z(19), FP_Z(18) => FP_Z(18)
                           , FP_Z(17) => FP_Z(17), FP_Z(16) => FP_Z(16), 
                           FP_Z(15) => FP_Z(15), FP_Z(14) => FP_Z(14), FP_Z(13)
                           => FP_Z(13), FP_Z(12) => FP_Z(12), FP_Z(11) => 
                           FP_Z(11), FP_Z(10) => FP_Z(10), FP_Z(9) => FP_Z(9), 
                           FP_Z(8) => FP_Z(8), FP_Z(7) => FP_Z(7), FP_Z(6) => 
                           FP_Z(6), FP_Z(5) => FP_Z(5), FP_Z(4) => FP_Z(4), 
                           FP_Z(3) => FP_Z(3), FP_Z(2) => FP_Z(2), FP_Z(1) => 
                           FP_Z(1), FP_Z(0) => FP_Z(0));
   MY_CLK_r_REG3_S4 : DFF_X1 port map( D => n8, CK => clk, Q => FP_Z(31), QN =>
                           n_2637);

end SYN_pipeline;
