library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

use IEEE.math_real.log2;
use IEEE.math_real.ceil;
use WORK.constants.all;


entity P4_ADDER is
		generic (	NBIT :	integer := NBIT;
					NBIT_PER_BLOCK: integer := NBIT_PER_BLOCK;
					NBLOCKS:	integer := NBLOCKS);
		port (	A 	:	in	std_logic_vector(NBIT-1 downto 0);
				B 	:	in	std_logic_vector(NBIT-1 downto 0);
				Cin :	in	std_logic;
				S 	:	out	std_logic_vector(NBIT-1 downto 0);
				Cout :	out	std_logic);
end P4_ADDER;


architecture STRUCTURAL of P4_ADDER is
-----------------------------COMPONENTS-------------------------------

component CARRY_GENERATOR 
		generic ( NBIT :		integer := NBIT;
				NBIT_PER_BLOCK: integer := NBIT_PER_BLOCK);
		port (
			A :		in	std_logic_vector(NBIT -1 downto 0);
			B :		in	std_logic_vector(NBIT -1 downto 0);
			Cin :	in	std_logic;
			Co :	out	std_logic_vector((NBIT/NBIT_PER_BLOCK) downto 0) );
end component;


component SUM_GENERATOR 
		generic (	NBIT_PER_BLOCK: integer := NBIT_PER_BLOCK;
					NBLOCKS:	integer := NBLOCKS); 
		port (	A:	in	std_logic_vector(NBIT_PER_BLOCK*NBLOCKS-1 downto 0);
				B:	in	std_logic_vector(NBIT_PER_BLOCK*NBLOCKS-1 downto 0);
				Ci:	in	std_logic_vector(NBLOCKS-1 downto 0);
				S:	out	std_logic_vector(NBIT_PER_BLOCK*NBLOCKS-1 downto 0));
end component;

-----------------------------END COMPONENTS---------------------------

-------------------------------SIGNALS--------------------------------

signal carry_out :std_logic_vector (NBLOCKS downto 0 ); --NBLOCK +1 to take into account also Cin=C0



-----------------------------END SIGNALS-------------------------------



begin

	CARRY_GEN_INST: CARRY_GENERATOR generic map (NBIT_PER_BLOCK => NBIT_PER_BLOCK, NBIT => NBIT_PER_BLOCK*NBLOCKS ) --defined in constants
									port map	(	A => A, 
													B => B,
													Cin => Cin,
													Co => carry_out);

	SUM_GEN_INST : SUM_GENERATOR 	generic map (NBIT_PER_BLOCK => NBIT_PER_BLOCK, NBLOCKS =>NBLOCKS)
								 	port map	(	A => A,
													B => B,
													Ci => carry_out (NBLOCKS -1 downto 0),
													S => S	);


	Cout <= carry_out (NBLOCKS); --final carry out is generated by carry_generator and it is the MSB of the signal connecting the SUM and CARRY GENERATORS



end STRUCTURAL;
