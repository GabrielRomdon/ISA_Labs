package CONSTANTS is
   constant NBIT_PER_BLOCK : integer := 2;
   constant NBLOCKS : integer := 32;
   constant NBIT : integer := NBLOCKS*NBIT_PER_BLOCK;
end CONSTANTS;
