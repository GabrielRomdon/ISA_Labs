
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_FPmul is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_FPmul;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPround_SIG_width28_DW01_inc_1 is

   port( A : in std_logic_vector (24 downto 0);  SUM : out std_logic_vector (24
         downto 0));

end FPround_SIG_width28_DW01_inc_1;

architecture SYN_USE_DEFA_ARCH_NAME of FPround_SIG_width28_DW01_inc_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n6, n7, n11, n14, n15, n16, n17, n18, n19, n23, n26, n27, n28
      , n29, n31, n35, n38, n39, n40, n41, n50, n51, n52, n56, n57, n61, n62, 
      n63, n68, n71, n72, n73, n74, n76, n80, n83, n84, n85, n86, n94, n95, n96
      , n97, n101, n105, n106, n113, n114, n115, n116, n122, n123, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194 : 
      std_logic;

begin
   
   U154 : AND2_X1 port map( A1 => n28, A2 => n6, ZN => n181);
   U155 : XNOR2_X1 port map( A => n182, B => A(3), ZN => SUM(3));
   U156 : NAND2_X1 port map( A1 => n122, A2 => A(2), ZN => n182);
   U157 : XOR2_X1 port map( A => n183, B => A(5), Z => SUM(5));
   U158 : NOR2_X1 port map( A1 => n114, A2 => n113, ZN => n183);
   U159 : XOR2_X1 port map( A => n184, B => A(6), Z => SUM(6));
   U160 : NOR2_X1 port map( A1 => n114, A2 => n105, ZN => n184);
   U161 : XOR2_X1 port map( A => n185, B => A(7), Z => SUM(7));
   U162 : NOR2_X1 port map( A1 => n114, A2 => n101, ZN => n185);
   U163 : XNOR2_X1 port map( A => n186, B => A(9), ZN => SUM(9));
   U164 : NAND2_X1 port map( A1 => n94, A2 => A(8), ZN => n186);
   U165 : XNOR2_X1 port map( A => n187, B => A(11), ZN => SUM(11));
   U166 : NAND2_X1 port map( A1 => n94, A2 => n80, ZN => n187);
   U167 : XNOR2_X1 port map( A => n188, B => A(13), ZN => SUM(13));
   U168 : NAND2_X1 port map( A1 => n68, A2 => n94, ZN => n188);
   U169 : XNOR2_X1 port map( A => n189, B => A(14), ZN => SUM(14));
   U170 : NAND2_X1 port map( A1 => n61, A2 => n94, ZN => n189);
   U171 : XNOR2_X1 port map( A => n190, B => A(15), ZN => SUM(15));
   U172 : NAND2_X1 port map( A1 => n56, A2 => n94, ZN => n190);
   U173 : XNOR2_X1 port map( A => n191, B => A(17), ZN => SUM(17));
   U174 : NAND2_X1 port map( A1 => n1, A2 => A(16), ZN => n191);
   U175 : XNOR2_X1 port map( A => n192, B => A(19), ZN => SUM(19));
   U176 : NAND2_X1 port map( A1 => n1, A2 => n35, ZN => n192);
   U177 : XNOR2_X1 port map( A => n193, B => A(21), ZN => SUM(21));
   U178 : NAND2_X1 port map( A1 => n1, A2 => n23, ZN => n193);
   U179 : XNOR2_X1 port map( A => n194, B => A(23), ZN => SUM(23));
   U180 : NAND2_X1 port map( A1 => n11, A2 => n1, ZN => n194);
   U181 : INV_X1 port map( A => n95, ZN => n94);
   U182 : INV_X1 port map( A => n115, ZN => n114);
   U183 : INV_X1 port map( A => n73, ZN => n74);
   U184 : NAND2_X1 port map( A1 => n1, A2 => n181, ZN => n3);
   U185 : NOR2_X1 port map( A1 => n19, A2 => n7, ZN => n6);
   U186 : NOR2_X1 port map( A1 => n41, A2 => n38, ZN => n35);
   U187 : NOR2_X1 port map( A1 => n86, A2 => n83, ZN => n80);
   U188 : NOR2_X1 port map( A1 => n29, A2 => n26, ZN => n23);
   U189 : INV_X1 port map( A => n28, ZN => n29);
   U190 : INV_X1 port map( A => n123, ZN => n122);
   U191 : NOR2_X1 port map( A1 => n74, A2 => n62, ZN => n61);
   U192 : NOR2_X1 port map( A1 => n74, A2 => n71, ZN => n68);
   U193 : NOR2_X1 port map( A1 => n17, A2 => n14, ZN => n11);
   U194 : NAND2_X1 port map( A1 => n28, A2 => n18, ZN => n17);
   U195 : INV_X1 port map( A => n19, ZN => n18);
   U196 : NOR2_X1 port map( A1 => n50, A2 => n95, ZN => n1);
   U197 : NAND2_X1 port map( A1 => n73, A2 => n51, ZN => n50);
   U198 : NOR2_X1 port map( A1 => n62, A2 => n52, ZN => n51);
   U199 : NAND2_X1 port map( A1 => A(14), A2 => A(15), ZN => n52);
   U200 : NOR2_X1 port map( A1 => n41, A2 => n31, ZN => n28);
   U201 : NAND2_X1 port map( A1 => A(18), A2 => A(19), ZN => n31);
   U202 : NOR2_X1 port map( A1 => n86, A2 => n76, ZN => n73);
   U203 : NAND2_X1 port map( A1 => A(10), A2 => A(11), ZN => n76);
   U204 : NOR2_X1 port map( A1 => n116, A2 => n123, ZN => n115);
   U205 : NAND2_X1 port map( A1 => A(2), A2 => A(3), ZN => n116);
   U206 : XOR2_X1 port map( A => n1, B => A(16), Z => SUM(16));
   U207 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n41);
   U208 : NAND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n86);
   U209 : XOR2_X1 port map( A => n84, B => n83, Z => SUM(10));
   U210 : NAND2_X1 port map( A1 => n94, A2 => n85, ZN => n84);
   U211 : INV_X1 port map( A => n86, ZN => n85);
   U212 : XOR2_X1 port map( A => n72, B => n71, Z => SUM(12));
   U213 : NAND2_X1 port map( A1 => n94, A2 => n73, ZN => n72);
   U214 : XOR2_X1 port map( A => n39, B => n38, Z => SUM(18));
   U215 : NAND2_X1 port map( A1 => n1, A2 => n40, ZN => n39);
   U216 : INV_X1 port map( A => n41, ZN => n40);
   U217 : XOR2_X1 port map( A => n27, B => n26, Z => SUM(20));
   U218 : NAND2_X1 port map( A1 => n1, A2 => n28, ZN => n27);
   U219 : XOR2_X1 port map( A => n15, B => n14, Z => SUM(22));
   U220 : NAND2_X1 port map( A1 => n1, A2 => n16, ZN => n15);
   U221 : INV_X1 port map( A => n17, ZN => n16);
   U222 : INV_X1 port map( A => A(18), ZN => n38);
   U223 : INV_X1 port map( A => A(20), ZN => n26);
   U224 : INV_X1 port map( A => A(10), ZN => n83);
   U225 : INV_X1 port map( A => A(22), ZN => n14);
   U226 : INV_X1 port map( A => A(12), ZN => n71);
   U227 : INV_X1 port map( A => A(4), ZN => n113);
   U228 : XOR2_X1 port map( A => n114, B => n113, Z => SUM(4));
   U229 : NAND2_X1 port map( A1 => A(4), A2 => A(5), ZN => n105);
   U230 : NAND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n62);
   U231 : XOR2_X1 port map( A => n94, B => A(8), Z => SUM(8));
   U232 : NOR2_X1 port map( A1 => n74, A2 => n57, ZN => n56);
   U233 : NAND2_X1 port map( A1 => n63, A2 => A(14), ZN => n57);
   U234 : INV_X1 port map( A => n62, ZN => n63);
   U235 : NAND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n123);
   U236 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n19);
   U237 : NAND2_X1 port map( A1 => n106, A2 => A(6), ZN => n101);
   U238 : INV_X1 port map( A => n105, ZN => n106);
   U239 : NAND2_X1 port map( A1 => A(22), A2 => A(23), ZN => n7);
   U240 : NAND2_X1 port map( A1 => n96, A2 => n115, ZN => n95);
   U241 : NOR2_X1 port map( A1 => n105, A2 => n97, ZN => n96);
   U242 : NAND2_X1 port map( A1 => A(6), A2 => A(7), ZN => n97);
   U243 : XOR2_X1 port map( A => n122, B => A(2), Z => SUM(2));
   U244 : INV_X1 port map( A => A(0), ZN => SUM(0));
   U245 : XOR2_X1 port map( A => A(1), B => A(0), Z => SUM(1));
   U246 : XNOR2_X1 port map( A => n3, B => A(24), ZN => SUM(24));

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage2_DW01_add_0 is

   port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (7 downto 0);  CO : out std_logic);

end FPmul_stage2_DW01_add_0;

architecture SYN_rpl of FPmul_stage2_DW01_add_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n_1002 : std_logic;

begin
   
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           n_1002, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1 : OR2_X1 port map( A1 => B(0), A2 => A(0), ZN => carry_1_port);
   U2 : XNOR2_X1 port map( A => B(0), B => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_15;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n13, ZN => Y(3));
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U4 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U5 : INV_X1 port map( A => SEL, ZN => n5);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_14;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n13, ZN => Y(3));
   U2 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U3 : INV_X1 port map( A => SEL, ZN => n5);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_13;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n13, ZN => Y(3));
   U2 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U3 : INV_X1 port map( A => SEL, ZN => n5);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_12;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n13, ZN => Y(3));
   U2 : INV_X1 port map( A => n12, ZN => Y(2));
   U3 : INV_X1 port map( A => n11, ZN => Y(1));
   U4 : INV_X1 port map( A => n10, ZN => Y(0));
   U5 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U6 : INV_X1 port map( A => SEL, ZN => n5);
   U7 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U8 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_11;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_10;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_9;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_8;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_7;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_6;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_5;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_4;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_3;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_2;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_1;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : INV_X1 port map( A => SEL, ZN => n5);
   U2 : INV_X1 port map( A => n13, ZN => Y(3));
   U3 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n13);
   U4 : INV_X1 port map( A => n12, ZN => Y(2));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n12);
   U6 : INV_X1 port map( A => n11, ZN => Y(1));
   U7 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n11);
   U8 : INV_X1 port map( A => n10, ZN => Y(0));
   U9 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_31;

architecture SYN_STRUCTURAL of RCA_generic_N4_31 is

   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_124 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_123 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_122 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_121 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_30;

architecture SYN_STRUCTURAL of RCA_generic_N4_30 is

   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_120 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_119 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_118 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_117 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_29;

architecture SYN_STRUCTURAL of RCA_generic_N4_29 is

   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_116 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_115 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_114 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_113 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_28;

architecture SYN_STRUCTURAL of RCA_generic_N4_28 is

   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_112 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_111 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_110 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_109 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_27;

architecture SYN_STRUCTURAL of RCA_generic_N4_27 is

   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_108 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_107 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_106 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_105 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_26;

architecture SYN_STRUCTURAL of RCA_generic_N4_26 is

   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_104 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_103 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_102 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_101 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_25;

architecture SYN_STRUCTURAL of RCA_generic_N4_25 is

   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_100 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_99 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_98 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_97 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_24;

architecture SYN_STRUCTURAL of RCA_generic_N4_24 is

   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_96 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_95 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_94 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_93 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_23;

architecture SYN_STRUCTURAL of RCA_generic_N4_23 is

   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_92 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_91 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_90 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_89 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_22;

architecture SYN_STRUCTURAL of RCA_generic_N4_22 is

   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_88 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_87 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_86 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_85 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_21;

architecture SYN_STRUCTURAL of RCA_generic_N4_21 is

   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_84 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_83 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_82 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_81 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_20;

architecture SYN_STRUCTURAL of RCA_generic_N4_20 is

   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_80 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_79 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_78 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_77 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_19;

architecture SYN_STRUCTURAL of RCA_generic_N4_19 is

   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_76 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_75 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_74 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_73 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_18;

architecture SYN_STRUCTURAL of RCA_generic_N4_18 is

   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_72 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_71 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_70 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_69 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_17;

architecture SYN_STRUCTURAL of RCA_generic_N4_17 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_68 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_67 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_66 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_65 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_16;

architecture SYN_STRUCTURAL of RCA_generic_N4_16 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_15;

architecture SYN_STRUCTURAL of RCA_generic_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_14;

architecture SYN_STRUCTURAL of RCA_generic_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_13;

architecture SYN_STRUCTURAL of RCA_generic_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_12;

architecture SYN_STRUCTURAL of RCA_generic_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_11;

architecture SYN_STRUCTURAL of RCA_generic_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_10;

architecture SYN_STRUCTURAL of RCA_generic_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_9;

architecture SYN_STRUCTURAL of RCA_generic_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_8;

architecture SYN_STRUCTURAL of RCA_generic_N4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_7;

architecture SYN_STRUCTURAL of RCA_generic_N4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_6;

architecture SYN_STRUCTURAL of RCA_generic_N4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_5;

architecture SYN_STRUCTURAL of RCA_generic_N4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_4;

architecture SYN_STRUCTURAL of RCA_generic_N4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_3;

architecture SYN_STRUCTURAL of RCA_generic_N4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_2;

architecture SYN_STRUCTURAL of RCA_generic_N4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_1;

architecture SYN_STRUCTURAL of RCA_generic_N4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_15;

architecture SYN_STRUCTURAL of carry_select_N4_15 is

   component MUX21_GENERIC_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1003, n_1004 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_30 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1003);
   ADDER1 : RCA_generic_N4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1004);
   MUX : MUX21_GENERIC_N4_15 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_14;

architecture SYN_STRUCTURAL of carry_select_N4_14 is

   component MUX21_GENERIC_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1005, n_1006 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1005);
   ADDER1 : RCA_generic_N4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1006);
   MUX : MUX21_GENERIC_N4_14 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_13;

architecture SYN_STRUCTURAL of carry_select_N4_13 is

   component MUX21_GENERIC_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1007, n_1008 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1007);
   ADDER1 : RCA_generic_N4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1008);
   MUX : MUX21_GENERIC_N4_13 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_12;

architecture SYN_STRUCTURAL of carry_select_N4_12 is

   component MUX21_GENERIC_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1009, n_1010 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1009);
   ADDER1 : RCA_generic_N4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1010);
   MUX : MUX21_GENERIC_N4_12 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_11;

architecture SYN_STRUCTURAL of carry_select_N4_11 is

   component MUX21_GENERIC_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1011, n_1012 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1011);
   ADDER1 : RCA_generic_N4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1012);
   MUX : MUX21_GENERIC_N4_11 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_10;

architecture SYN_STRUCTURAL of carry_select_N4_10 is

   component MUX21_GENERIC_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1013, n_1014 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1013);
   ADDER1 : RCA_generic_N4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1014);
   MUX : MUX21_GENERIC_N4_10 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_9;

architecture SYN_STRUCTURAL of carry_select_N4_9 is

   component MUX21_GENERIC_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1015, n_1016 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1015);
   ADDER1 : RCA_generic_N4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1016);
   MUX : MUX21_GENERIC_N4_9 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_8;

architecture SYN_STRUCTURAL of carry_select_N4_8 is

   component MUX21_GENERIC_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1017, n_1018 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1017);
   ADDER1 : RCA_generic_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1018);
   MUX : MUX21_GENERIC_N4_8 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_7;

architecture SYN_STRUCTURAL of carry_select_N4_7 is

   component MUX21_GENERIC_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1019, n_1020 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1019);
   ADDER1 : RCA_generic_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1020);
   MUX : MUX21_GENERIC_N4_7 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_6;

architecture SYN_STRUCTURAL of carry_select_N4_6 is

   component MUX21_GENERIC_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1021, n_1022 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1021);
   ADDER1 : RCA_generic_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1022);
   MUX : MUX21_GENERIC_N4_6 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_5;

architecture SYN_STRUCTURAL of carry_select_N4_5 is

   component MUX21_GENERIC_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1023, n_1024 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1023);
   ADDER1 : RCA_generic_N4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1024);
   MUX : MUX21_GENERIC_N4_5 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_4;

architecture SYN_STRUCTURAL of carry_select_N4_4 is

   component MUX21_GENERIC_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1025, n_1026 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1025);
   ADDER1 : RCA_generic_N4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1026);
   MUX : MUX21_GENERIC_N4_4 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_3;

architecture SYN_STRUCTURAL of carry_select_N4_3 is

   component MUX21_GENERIC_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1027, n_1028 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1027);
   ADDER1 : RCA_generic_N4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1028);
   MUX : MUX21_GENERIC_N4_3 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_2;

architecture SYN_STRUCTURAL of carry_select_N4_2 is

   component MUX21_GENERIC_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1029, n_1030 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1029);
   ADDER1 : RCA_generic_N4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1030);
   MUX : MUX21_GENERIC_N4_2 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_1;

architecture SYN_STRUCTURAL of carry_select_N4_1 is

   component MUX21_GENERIC_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1031, n_1032 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1031);
   ADDER1 : RCA_generic_N4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1032);
   MUX : MUX21_GENERIC_N4_1 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_62 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_62;

architecture SYN_BEHAVIORAL of PG_GENERAL_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_61 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_61;

architecture SYN_BEHAVIORAL of PG_GENERAL_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_60 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_60;

architecture SYN_BEHAVIORAL of PG_GENERAL_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_59 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_59;

architecture SYN_BEHAVIORAL of PG_GENERAL_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_58 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_58;

architecture SYN_BEHAVIORAL of PG_GENERAL_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_57 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_57;

architecture SYN_BEHAVIORAL of PG_GENERAL_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_56 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_56;

architecture SYN_BEHAVIORAL of PG_GENERAL_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_55 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_55;

architecture SYN_BEHAVIORAL of PG_GENERAL_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_54 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_54;

architecture SYN_BEHAVIORAL of PG_GENERAL_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : OAI22_X1 port map( A1 => PG_ik(0), A2 => PG_ik(1), B1 => PG_k_1j(1), B2
                           => PG_ik(1), ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_53 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_53;

architecture SYN_BEHAVIORAL of PG_GENERAL_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_52 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_52;

architecture SYN_BEHAVIORAL of PG_GENERAL_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => PG_ik(0), Z => n1);
   U2 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => n1, ZN => PG_ij(0));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n2);
   U4 : INV_X1 port map( A => n2, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_51 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_51;

architecture SYN_BEHAVIORAL of PG_GENERAL_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_50 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_50;

architecture SYN_BEHAVIORAL of PG_GENERAL_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net39810, n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : OAI21_X1 port map( B1 => net39810, B2 => n1, A => n2, ZN => PG_ij(1));
   U3 : INV_X1 port map( A => PG_ik(0), ZN => net39810);
   U4 : INV_X1 port map( A => PG_k_1j(1), ZN => n1);
   U5 : INV_X1 port map( A => PG_ik(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_49 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_49;

architecture SYN_BEHAVIORAL of PG_GENERAL_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_48 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_48;

architecture SYN_BEHAVIORAL of PG_GENERAL_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => PG_ik(0), Z => n1);
   U2 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => n1, ZN => PG_ij(0));
   U3 : OAI22_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(1), B1 => PG_ik(0), B2
                           => PG_ik(1), ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_47 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_47;

architecture SYN_BEHAVIORAL of PG_GENERAL_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_46 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_46;

architecture SYN_BEHAVIORAL of PG_GENERAL_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PG_ij(1));
   U2 : INV_X1 port map( A => PG_ik(0), ZN => n1);
   U3 : INV_X1 port map( A => PG_k_1j(1), ZN => n2);
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n3);
   U5 : CLKBUF_X1 port map( A => PG_ik(0), Z => n4);
   U6 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => n4, ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_45 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_45;

architecture SYN_BEHAVIORAL of PG_GENERAL_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PG_ij(1));
   U2 : INV_X1 port map( A => PG_ik(0), ZN => n1);
   U3 : INV_X1 port map( A => PG_k_1j(1), ZN => n2);
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n3);
   U5 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_44 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_44;

architecture SYN_BEHAVIORAL of PG_GENERAL_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_43 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_43;

architecture SYN_BEHAVIORAL of PG_GENERAL_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_42 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_42;

architecture SYN_BEHAVIORAL of PG_GENERAL_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_41 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_41;

architecture SYN_BEHAVIORAL of PG_GENERAL_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_40 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_40;

architecture SYN_BEHAVIORAL of PG_GENERAL_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_39 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_39;

architecture SYN_BEHAVIORAL of PG_GENERAL_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_38 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_38;

architecture SYN_BEHAVIORAL of PG_GENERAL_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_37 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_37;

architecture SYN_BEHAVIORAL of PG_GENERAL_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_36 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_36;

architecture SYN_BEHAVIORAL of PG_GENERAL_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U2 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U3 : INV_X1 port map( A => n3, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_35 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_35;

architecture SYN_BEHAVIORAL of PG_GENERAL_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_34 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_34;

architecture SYN_BEHAVIORAL of PG_GENERAL_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U2 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U3 : INV_X1 port map( A => n3, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_33 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_33;

architecture SYN_BEHAVIORAL of PG_GENERAL_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_32 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_32;

architecture SYN_BEHAVIORAL of PG_GENERAL_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_31 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_31;

architecture SYN_BEHAVIORAL of PG_GENERAL_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_30 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_30;

architecture SYN_BEHAVIORAL of PG_GENERAL_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_29 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_29;

architecture SYN_BEHAVIORAL of PG_GENERAL_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_28 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_28;

architecture SYN_BEHAVIORAL of PG_GENERAL_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n2, A2 => PG_ik(1), ZN => PG_ij(1));
   U2 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n2);
   U3 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_27 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_27;

architecture SYN_BEHAVIORAL of PG_GENERAL_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PG_ij(1));
   U2 : INV_X1 port map( A => PG_k_1j(1), ZN => n1);
   U3 : INV_X1 port map( A => PG_ik(0), ZN => n2);
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n3);
   U5 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_26 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_26;

architecture SYN_BEHAVIORAL of PG_GENERAL_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net39840, n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : OAI21_X1 port map( B1 => n1, B2 => net39840, A => n2, ZN => PG_ij(1));
   U3 : INV_X1 port map( A => PG_k_1j(1), ZN => n1);
   U4 : INV_X1 port map( A => PG_ik(0), ZN => net39840);
   U5 : INV_X1 port map( A => PG_ik(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_25 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_25;

architecture SYN_BEHAVIORAL of PG_GENERAL_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_24 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_24;

architecture SYN_BEHAVIORAL of PG_GENERAL_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_23 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_23;

architecture SYN_BEHAVIORAL of PG_GENERAL_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_22 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_22;

architecture SYN_BEHAVIORAL of PG_GENERAL_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_21 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_21;

architecture SYN_BEHAVIORAL of PG_GENERAL_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_20 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_20;

architecture SYN_BEHAVIORAL of PG_GENERAL_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_19 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_19;

architecture SYN_BEHAVIORAL of PG_GENERAL_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_18 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_18;

architecture SYN_BEHAVIORAL of PG_GENERAL_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_17 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_17;

architecture SYN_BEHAVIORAL of PG_GENERAL_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_16 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_16;

architecture SYN_BEHAVIORAL of PG_GENERAL_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : OR2_X2 port map( A1 => n2, A2 => PG_ik(1), ZN => PG_ij(1));
   U2 : AND2_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(0), ZN => n2);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_15 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_15;

architecture SYN_BEHAVIORAL of PG_GENERAL_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n1, A2 => PG_ik(1), ZN => PG_ij(1));
   U2 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n1);
   U3 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_14 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_14;

architecture SYN_BEHAVIORAL of PG_GENERAL_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_13 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_13;

architecture SYN_BEHAVIORAL of PG_GENERAL_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_12 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_12;

architecture SYN_BEHAVIORAL of PG_GENERAL_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_11 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_11;

architecture SYN_BEHAVIORAL of PG_GENERAL_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_10 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_10;

architecture SYN_BEHAVIORAL of PG_GENERAL_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_9 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_9;

architecture SYN_BEHAVIORAL of PG_GENERAL_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_8 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_8;

architecture SYN_BEHAVIORAL of PG_GENERAL_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U2 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_7 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_7;

architecture SYN_BEHAVIORAL of PG_GENERAL_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_6 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_6;

architecture SYN_BEHAVIORAL of PG_GENERAL_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_5 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_5;

architecture SYN_BEHAVIORAL of PG_GENERAL_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_4 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_4;

architecture SYN_BEHAVIORAL of PG_GENERAL_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_3 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_3;

architecture SYN_BEHAVIORAL of PG_GENERAL_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_2 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_2;

architecture SYN_BEHAVIORAL of PG_GENERAL_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);
   U2 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_1 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_1;

architecture SYN_BEHAVIORAL of PG_GENERAL_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_ij(1));
   U2 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U3 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_16 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_16;

architecture SYN_BEHAVIORAL of G_GENERAL_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_15 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_15;

architecture SYN_BEHAVIORAL of G_GENERAL_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_14 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_14;

architecture SYN_BEHAVIORAL of G_GENERAL_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => G_k_1j, A => PG_ik(1), ZN => 
                           n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_13 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_13;

architecture SYN_BEHAVIORAL of G_GENERAL_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_12 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_12;

architecture SYN_BEHAVIORAL of G_GENERAL_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_11 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_11;

architecture SYN_BEHAVIORAL of G_GENERAL_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_10 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_10;

architecture SYN_BEHAVIORAL of G_GENERAL_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_9 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_9;

architecture SYN_BEHAVIORAL of G_GENERAL_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OR2_X2 port map( A1 => PG_ik(1), A2 => n1, ZN => G_ij);
   U2 : AND2_X1 port map( A1 => G_k_1j, A2 => PG_ik(0), ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_8 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_8;

architecture SYN_BEHAVIORAL of G_GENERAL_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_7 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_7;

architecture SYN_BEHAVIORAL of G_GENERAL_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_6 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_6;

architecture SYN_BEHAVIORAL of G_GENERAL_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_5 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_5;

architecture SYN_BEHAVIORAL of G_GENERAL_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => G_k_1j, A => PG_ik(1), ZN => 
                           n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_4 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_4;

architecture SYN_BEHAVIORAL of G_GENERAL_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => G_k_1j, A => PG_ik(1), ZN => 
                           n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_3 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_3;

architecture SYN_BEHAVIORAL of G_GENERAL_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => G_k_1j, A => PG_ik(1), ZN => 
                           n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_2 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_2;

architecture SYN_BEHAVIORAL of G_GENERAL_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => G_k_1j, A => PG_ik(1), ZN => 
                           n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_1 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_1;

architecture SYN_BEHAVIORAL of G_GENERAL_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => G_k_1j, A => PG_ik(1), ZN => 
                           n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_63 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_63;

architecture SYN_BEHAVIORAL of PG_NET_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_62 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_62;

architecture SYN_BEHAVIORAL of PG_NET_62 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_61 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_61;

architecture SYN_BEHAVIORAL of PG_NET_61 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_60 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_60;

architecture SYN_BEHAVIORAL of PG_NET_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_59 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_59;

architecture SYN_BEHAVIORAL of PG_NET_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_58 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_58;

architecture SYN_BEHAVIORAL of PG_NET_58 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_57 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_57;

architecture SYN_BEHAVIORAL of PG_NET_57 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_56 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_56;

architecture SYN_BEHAVIORAL of PG_NET_56 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_55 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_55;

architecture SYN_BEHAVIORAL of PG_NET_55 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_54 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_54;

architecture SYN_BEHAVIORAL of PG_NET_54 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_53 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_53;

architecture SYN_BEHAVIORAL of PG_NET_53 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_52 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_52;

architecture SYN_BEHAVIORAL of PG_NET_52 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_51 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_51;

architecture SYN_BEHAVIORAL of PG_NET_51 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_50 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_50;

architecture SYN_BEHAVIORAL of PG_NET_50 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_49 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_49;

architecture SYN_BEHAVIORAL of PG_NET_49 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_48 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_48;

architecture SYN_BEHAVIORAL of PG_NET_48 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_47 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_47;

architecture SYN_BEHAVIORAL of PG_NET_47 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_46 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_46;

architecture SYN_BEHAVIORAL of PG_NET_46 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_45 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_45;

architecture SYN_BEHAVIORAL of PG_NET_45 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_44 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_44;

architecture SYN_BEHAVIORAL of PG_NET_44 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_43 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_43;

architecture SYN_BEHAVIORAL of PG_NET_43 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_42 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_42;

architecture SYN_BEHAVIORAL of PG_NET_42 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_41 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_41;

architecture SYN_BEHAVIORAL of PG_NET_41 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_40 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_40;

architecture SYN_BEHAVIORAL of PG_NET_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_39 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_39;

architecture SYN_BEHAVIORAL of PG_NET_39 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_38 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_38;

architecture SYN_BEHAVIORAL of PG_NET_38 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_37 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_37;

architecture SYN_BEHAVIORAL of PG_NET_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => B, ZN => n1);
   U2 : XNOR2_X1 port map( A => A, B => n1, ZN => P_OUT);
   U3 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_36 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_36;

architecture SYN_BEHAVIORAL of PG_NET_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_35 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_35;

architecture SYN_BEHAVIORAL of PG_NET_35 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net27182, net27183 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => net27182);
   U3 : INV_X1 port map( A => B, ZN => net27183);
   U4 : NOR2_X1 port map( A1 => net27182, A2 => net27183, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_34 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_34;

architecture SYN_BEHAVIORAL of PG_NET_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_33 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_33;

architecture SYN_BEHAVIORAL of PG_NET_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_32 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_32;

architecture SYN_BEHAVIORAL of PG_NET_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_31 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_31;

architecture SYN_BEHAVIORAL of PG_NET_31 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_30 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_30;

architecture SYN_BEHAVIORAL of PG_NET_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_29 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_29;

architecture SYN_BEHAVIORAL of PG_NET_29 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_28 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_28;

architecture SYN_BEHAVIORAL of PG_NET_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_27 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_27;

architecture SYN_BEHAVIORAL of PG_NET_27 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net27166, net27167 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => net27166);
   U3 : INV_X1 port map( A => B, ZN => net27167);
   U4 : NOR2_X1 port map( A1 => net27166, A2 => net27167, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_26 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_26;

architecture SYN_BEHAVIORAL of PG_NET_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_25 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_25;

architecture SYN_BEHAVIORAL of PG_NET_25 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_24 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_24;

architecture SYN_BEHAVIORAL of PG_NET_24 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_23 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_23;

architecture SYN_BEHAVIORAL of PG_NET_23 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_22 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_22;

architecture SYN_BEHAVIORAL of PG_NET_22 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n2, ZN => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_21 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_21;

architecture SYN_BEHAVIORAL of PG_NET_21 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n2, ZN => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_20 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_20;

architecture SYN_BEHAVIORAL of PG_NET_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_19 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_19;

architecture SYN_BEHAVIORAL of PG_NET_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_18 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_18;

architecture SYN_BEHAVIORAL of PG_NET_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_17 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_17;

architecture SYN_BEHAVIORAL of PG_NET_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_16 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_16;

architecture SYN_BEHAVIORAL of PG_NET_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_15 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_15;

architecture SYN_BEHAVIORAL of PG_NET_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_14 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_14;

architecture SYN_BEHAVIORAL of PG_NET_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_13 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_13;

architecture SYN_BEHAVIORAL of PG_NET_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_12 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_12;

architecture SYN_BEHAVIORAL of PG_NET_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_11 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_11;

architecture SYN_BEHAVIORAL of PG_NET_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_10 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_10;

architecture SYN_BEHAVIORAL of PG_NET_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_9 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_9;

architecture SYN_BEHAVIORAL of PG_NET_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_8 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_8;

architecture SYN_BEHAVIORAL of PG_NET_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_7 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_7;

architecture SYN_BEHAVIORAL of PG_NET_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_6 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_6;

architecture SYN_BEHAVIORAL of PG_NET_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_5 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_5;

architecture SYN_BEHAVIORAL of PG_NET_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_4 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_4;

architecture SYN_BEHAVIORAL of PG_NET_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_3 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_3;

architecture SYN_BEHAVIORAL of PG_NET_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_2 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_2;

architecture SYN_BEHAVIORAL of PG_NET_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_1 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_1;

architecture SYN_BEHAVIORAL of PG_NET_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_607 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_607;

architecture SYN_BEHAVIORAL of FA_607 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net29057, net29058, net29059, net29060, n1, n2, n3, n4, n5 : 
      std_logic;

begin
   
   U1 : BUF_X1 port map( A => B, Z => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U3 : NAND2_X1 port map( A1 => net29057, A2 => net29058, ZN => n2);
   U4 : NAND2_X1 port map( A1 => net29059, A2 => net29060, ZN => n3);
   U5 : AND2_X2 port map( A1 => n3, A2 => n2, ZN => Co);
   U6 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U7 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U8 : INV_X1 port map( A => A, ZN => net29057);
   U9 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => net29059);
   U10 : INV_X1 port map( A => n4, ZN => net29058);
   U11 : INV_X1 port map( A => n1, ZN => net29060);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_606 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_606;

architecture SYN_BEHAVIORAL of FA_606 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n2);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n7);
   U4 : XNOR2_X1 port map( A => n7, B => A, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n6);
   U6 : INV_X1 port map( A => n1, ZN => n5);
   U7 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U8 : INV_X1 port map( A => n2, ZN => n3);
   U9 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_605 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_605;

architecture SYN_BEHAVIORAL of FA_605 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n3);
   U2 : INV_X1 port map( A => n3, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n2);
   U5 : AND2_X2 port map( A1 => n1, A2 => n2, ZN => Co);
   U6 : CLKBUF_X1 port map( A => B, Z => n4);
   U7 : XNOR2_X1 port map( A => n9, B => Ci, ZN => S);
   U8 : XNOR2_X1 port map( A => B, B => A, ZN => n9);
   U9 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n8);
   U10 : INV_X1 port map( A => Ci, ZN => n7);
   U11 : INV_X1 port map( A => n4, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_604 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_604;

architecture SYN_BEHAVIORAL of FA_604 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_603 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_603;

architecture SYN_BEHAVIORAL of FA_603 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29038, net29039, net29040, net34131, n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);
   U2 : BUF_X1 port map( A => B, Z => net34131);
   U3 : NAND2_X1 port map( A1 => n4, A2 => net29038, ZN => n1);
   U4 : NAND2_X1 port map( A1 => net29039, A2 => net29040, ZN => n2);
   U5 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U7 : INV_X1 port map( A => Ci, ZN => net29038);
   U8 : INV_X1 port map( A => A, ZN => net29039);
   U9 : NAND2_X1 port map( A1 => net34131, A2 => A, ZN => n4);
   U10 : INV_X1 port map( A => net34131, ZN => net29040);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_602 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_602;

architecture SYN_BEHAVIORAL of FA_602 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n2);
   U3 : AND2_X2 port map( A1 => n1, A2 => n2, ZN => Co);
   U4 : XNOR2_X1 port map( A => B, B => n7, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n5);
   U8 : INV_X1 port map( A => A, ZN => n4);
   U9 : INV_X1 port map( A => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_601 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_601;

architecture SYN_BEHAVIORAL of FA_601 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_600 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_600;

architecture SYN_BEHAVIORAL of FA_600 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_599 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_599;

architecture SYN_BEHAVIORAL of FA_599 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_598 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_598;

architecture SYN_BEHAVIORAL of FA_598 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n_1033 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : INV_X1 port map( A => B, ZN => n2);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U5 : FA_X1 port map( A => Ci, B => A, CI => B, CO => n_1033, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_597 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_597;

architecture SYN_BEHAVIORAL of FA_597 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_596 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_596;

architecture SYN_BEHAVIORAL of FA_596 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI22_X2 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_595 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_595;

architecture SYN_BEHAVIORAL of FA_595 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_594 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_594;

architecture SYN_BEHAVIORAL of FA_594 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_593 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_593;

architecture SYN_BEHAVIORAL of FA_593 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_592 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_592;

architecture SYN_BEHAVIORAL of FA_592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n2, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : CLKBUF_X1 port map( A => B, Z => n2);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_591 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_591;

architecture SYN_BEHAVIORAL of FA_591 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28980, net28981, net28982, net28983, net34026, net34175, n1, n2, 
      n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : INV_X1 port map( A => B, ZN => net28981);
   U4 : CLKBUF_X1 port map( A => Ci, Z => net34026);
   U5 : INV_X1 port map( A => A, ZN => net28980);
   U6 : NAND2_X1 port map( A1 => net34175, A2 => A, ZN => net28982);
   U7 : NAND2_X1 port map( A1 => net28980, A2 => net28981, ZN => n2);
   U8 : NAND2_X1 port map( A1 => net28982, A2 => net28983, ZN => n3);
   U9 : AND2_X2 port map( A1 => n2, A2 => n3, ZN => Co);
   U10 : INV_X1 port map( A => net28981, ZN => net34175);
   U11 : INV_X1 port map( A => net34026, ZN => net28983);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_590 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_590;

architecture SYN_BEHAVIORAL of FA_590 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n2, B2 => n3, A => n1, ZN => Co);
   U2 : INV_X1 port map( A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U5 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U6 : XOR2_X1 port map( A => Ci, B => n4, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_589 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_589;

architecture SYN_BEHAVIORAL of FA_589 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => A, ZN => n2);
   U7 : INV_X1 port map( A => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_588 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_588;

architecture SYN_BEHAVIORAL of FA_588 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_587 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_587;

architecture SYN_BEHAVIORAL of FA_587 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U4 : INV_X1 port map( A => n1, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_586 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_586;

architecture SYN_BEHAVIORAL of FA_586 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_585 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_585;

architecture SYN_BEHAVIORAL of FA_585 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_584 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_584;

architecture SYN_BEHAVIORAL of FA_584 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_583 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_583;

architecture SYN_BEHAVIORAL of FA_583 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => n1, B => n4, ZN => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_582 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_582;

architecture SYN_BEHAVIORAL of FA_582 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_581 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_581;

architecture SYN_BEHAVIORAL of FA_581 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_580 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_580;

architecture SYN_BEHAVIORAL of FA_580 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n1);
   U2 : XNOR2_X1 port map( A => n2, B => n1, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n2);
   U4 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => Co);
   U5 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_579 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_579;

architecture SYN_BEHAVIORAL of FA_579 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n2, ZN => S);
   U3 : XNOR2_X1 port map( A => n1, B => B, ZN => n2);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U5 : AND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => Ci, B2 => n3, ZN => n5);
   U7 : INV_X1 port map( A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_578 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_578;

architecture SYN_BEHAVIORAL of FA_578 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_577 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_577;

architecture SYN_BEHAVIORAL of FA_577 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_576 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_576;

architecture SYN_BEHAVIORAL of FA_576 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_575 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_575;

architecture SYN_BEHAVIORAL of FA_575 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_574 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_574;

architecture SYN_BEHAVIORAL of FA_574 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_573 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_573;

architecture SYN_BEHAVIORAL of FA_573 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U3 : AOI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_572 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_572;

architecture SYN_BEHAVIORAL of FA_572 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_571 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_571;

architecture SYN_BEHAVIORAL of FA_571 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : CLKBUF_X1 port map( A => B, Z => n2);
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => n1, ZN => n5);
   U6 : INV_X1 port map( A => n2, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n2, B2 => n1, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_570 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_570;

architecture SYN_BEHAVIORAL of FA_570 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : CLKBUF_X1 port map( A => B, Z => n2);
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => n1, ZN => n5);
   U6 : INV_X1 port map( A => n2, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n2, B2 => n1, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_569 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_569;

architecture SYN_BEHAVIORAL of FA_569 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_568 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_568;

architecture SYN_BEHAVIORAL of FA_568 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_567 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_567;

architecture SYN_BEHAVIORAL of FA_567 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_566 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_566;

architecture SYN_BEHAVIORAL of FA_566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_565 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_565;

architecture SYN_BEHAVIORAL of FA_565 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_564 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_564;

architecture SYN_BEHAVIORAL of FA_564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_563 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_563;

architecture SYN_BEHAVIORAL of FA_563 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_562 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_562;

architecture SYN_BEHAVIORAL of FA_562 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_561 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_561;

architecture SYN_BEHAVIORAL of FA_561 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_560 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_560;

architecture SYN_BEHAVIORAL of FA_560 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U4 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U5 : XNOR2_X1 port map( A => A, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_559 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_559;

architecture SYN_BEHAVIORAL of FA_559 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net28830, net28833, net28834, net34005, net34078, n1, n2, n3, n4, n5 
      : std_logic;

begin
   
   U1 : BUF_X1 port map( A => B, Z => n1);
   U2 : XNOR2_X1 port map( A => n2, B => n1, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U4 : NAND2_X1 port map( A1 => net34078, A2 => n1, ZN => net28830);
   U5 : INV_X1 port map( A => B, ZN => net28833);
   U6 : INV_X1 port map( A => A, ZN => net28834);
   U7 : BUF_X1 port map( A => Ci, Z => net34005);
   U8 : INV_X1 port map( A => net28834, ZN => net34078);
   U9 : NAND2_X1 port map( A1 => n5, A2 => net28830, ZN => Co);
   U10 : XNOR2_X1 port map( A => n4, B => n3, ZN => n5);
   U11 : NAND2_X1 port map( A1 => net34005, A2 => net28833, ZN => n3);
   U12 : NAND2_X1 port map( A1 => net34005, A2 => net28834, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_558 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_558;

architecture SYN_BEHAVIORAL of FA_558 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => n1);
   U2 : CLKBUF_X1 port map( A => A, Z => n2);
   U3 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U5 : INV_X1 port map( A => n2, ZN => n6);
   U6 : INV_X1 port map( A => B, ZN => n5);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => n4);
   U8 : INV_X1 port map( A => Ci, ZN => n3);
   U9 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_557 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_557;

architecture SYN_BEHAVIORAL of FA_557 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28819, net28820, net28821, net28822, net34181, net34316, n1 : 
      std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => net28821);
   U4 : CLKBUF_X1 port map( A => Ci, Z => net34316);
   U5 : NAND2_X1 port map( A1 => B, A2 => net34181, ZN => net28819);
   U6 : INV_X1 port map( A => B, ZN => net28822);
   U7 : INV_X1 port map( A => net28821, ZN => net34181);
   U8 : INV_X1 port map( A => net34316, ZN => net28820);
   U9 : AOI22_X1 port map( A1 => net28819, A2 => net28820, B1 => net28821, B2 
                           => net28822, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_556 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_556;

architecture SYN_BEHAVIORAL of FA_556 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : AOI22_X2 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => n1, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : NAND2_X1 port map( A1 => B, A2 => n1, ZN => n3);
   U8 : INV_X1 port map( A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_555 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_555;

architecture SYN_BEHAVIORAL of FA_555 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net28809, net28810, net28811, net28812, net31437, n1 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => A, Z => net31437);
   U2 : AOI22_X2 port map( A1 => net28809, A2 => net28810, B1 => net28811, B2 
                           => net28812, ZN => Co);
   U3 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U5 : NAND2_X1 port map( A1 => B, A2 => net31437, ZN => net28809);
   U6 : INV_X1 port map( A => B, ZN => net28812);
   U7 : INV_X1 port map( A => Ci, ZN => net28810);
   U8 : INV_X1 port map( A => net31437, ZN => net28811);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_554 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_554;

architecture SYN_BEHAVIORAL of FA_554 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : INV_X1 port map( A => n5, ZN => n2);
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n1, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n1, B2 => n2, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_553 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_553;

architecture SYN_BEHAVIORAL of FA_553 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n1);
   U2 : XNOR2_X1 port map( A => n8, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n8);
   U4 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U6 : XNOR2_X1 port map( A => n5, B => n4, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => n5);
   U8 : NAND2_X1 port map( A1 => n1, A2 => n3, ZN => n4);
   U9 : INV_X1 port map( A => A, ZN => n2);
   U10 : INV_X1 port map( A => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_552 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_552;

architecture SYN_BEHAVIORAL of FA_552 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_551 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_551;

architecture SYN_BEHAVIORAL of FA_551 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_550 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_550;

architecture SYN_BEHAVIORAL of FA_550 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_549 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_549;

architecture SYN_BEHAVIORAL of FA_549 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : XNOR2_X1 port map( A => n1, B => n4, ZN => S);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_548 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_548;

architecture SYN_BEHAVIORAL of FA_548 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_547 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_547;

architecture SYN_BEHAVIORAL of FA_547 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => n1, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_546 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_546;

architecture SYN_BEHAVIORAL of FA_546 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_545 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_545;

architecture SYN_BEHAVIORAL of FA_545 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_544 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_544;

architecture SYN_BEHAVIORAL of FA_544 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_543 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_543;

architecture SYN_BEHAVIORAL of FA_543 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_542 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_542;

architecture SYN_BEHAVIORAL of FA_542 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_541 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_541;

architecture SYN_BEHAVIORAL of FA_541 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_540 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_540;

architecture SYN_BEHAVIORAL of FA_540 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_539 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_539;

architecture SYN_BEHAVIORAL of FA_539 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_538 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_538;

architecture SYN_BEHAVIORAL of FA_538 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_537 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_537;

architecture SYN_BEHAVIORAL of FA_537 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_536 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_536;

architecture SYN_BEHAVIORAL of FA_536 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_535 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_535;

architecture SYN_BEHAVIORAL of FA_535 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_534 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_534;

architecture SYN_BEHAVIORAL of FA_534 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_533 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_533;

architecture SYN_BEHAVIORAL of FA_533 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_532 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_532;

architecture SYN_BEHAVIORAL of FA_532 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_531 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_531;

architecture SYN_BEHAVIORAL of FA_531 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_530 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_530;

architecture SYN_BEHAVIORAL of FA_530 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_529 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_529;

architecture SYN_BEHAVIORAL of FA_529 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_528 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_528;

architecture SYN_BEHAVIORAL of FA_528 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_527 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_527;

architecture SYN_BEHAVIORAL of FA_527 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U2 : CLKBUF_X1 port map( A => A, Z => n2);
   U3 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U5 : INV_X1 port map( A => n2, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => n2, A => n1, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_526 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_526;

architecture SYN_BEHAVIORAL of FA_526 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => B, Z => n1);
   U2 : XNOR2_X1 port map( A => n2, B => n1, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_525 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_525;

architecture SYN_BEHAVIORAL of FA_525 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n2);
   U3 : XNOR2_X1 port map( A => n7, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => A, ZN => n7);
   U5 : NAND2_X1 port map( A1 => B, A2 => n1, ZN => n6);
   U6 : INV_X1 port map( A => n2, ZN => n5);
   U7 : INV_X1 port map( A => A, ZN => n4);
   U8 : INV_X1 port map( A => B, ZN => n3);
   U9 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_524 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_524;

architecture SYN_BEHAVIORAL of FA_524 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n2);
   U3 : XNOR2_X1 port map( A => n7, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => A, ZN => n7);
   U5 : NAND2_X1 port map( A1 => B, A2 => n1, ZN => n6);
   U6 : INV_X1 port map( A => n2, ZN => n5);
   U7 : INV_X1 port map( A => A, ZN => n4);
   U8 : INV_X1 port map( A => B, ZN => n3);
   U9 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_523 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_523;

architecture SYN_BEHAVIORAL of FA_523 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_522 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_522;

architecture SYN_BEHAVIORAL of FA_522 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_521 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_521;

architecture SYN_BEHAVIORAL of FA_521 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => n1, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n1, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_520 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_520;

architecture SYN_BEHAVIORAL of FA_520 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => n1);
   U2 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n1, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_519 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_519;

architecture SYN_BEHAVIORAL of FA_519 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_518 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_518;

architecture SYN_BEHAVIORAL of FA_518 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => n1);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => A, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_517 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_517;

architecture SYN_BEHAVIORAL of FA_517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_516 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_516;

architecture SYN_BEHAVIORAL of FA_516 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_515 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_515;

architecture SYN_BEHAVIORAL of FA_515 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_514 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_514;

architecture SYN_BEHAVIORAL of FA_514 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_513 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_513;

architecture SYN_BEHAVIORAL of FA_513 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_512 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_512;

architecture SYN_BEHAVIORAL of FA_512 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_511;

architecture SYN_BEHAVIORAL of FA_511 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_510;

architecture SYN_BEHAVIORAL of FA_510 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_509;

architecture SYN_BEHAVIORAL of FA_509 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_508;

architecture SYN_BEHAVIORAL of FA_508 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_507;

architecture SYN_BEHAVIORAL of FA_507 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_506;

architecture SYN_BEHAVIORAL of FA_506 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_505;

architecture SYN_BEHAVIORAL of FA_505 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_504;

architecture SYN_BEHAVIORAL of FA_504 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_503;

architecture SYN_BEHAVIORAL of FA_503 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_502;

architecture SYN_BEHAVIORAL of FA_502 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_501;

architecture SYN_BEHAVIORAL of FA_501 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_500;

architecture SYN_BEHAVIORAL of FA_500 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => B, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_499;

architecture SYN_BEHAVIORAL of FA_499 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_498;

architecture SYN_BEHAVIORAL of FA_498 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_497;

architecture SYN_BEHAVIORAL of FA_497 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_496;

architecture SYN_BEHAVIORAL of FA_496 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => n1, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n1, B2 => B, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_495;

architecture SYN_BEHAVIORAL of FA_495 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_494;

architecture SYN_BEHAVIORAL of FA_494 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28552, net28553, net28554, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net28554);
   U4 : INV_X1 port map( A => A, ZN => net28552);
   U5 : INV_X1 port map( A => B, ZN => net28553);
   U6 : OAI21_X1 port map( B1 => net28552, B2 => net28553, A => net28554, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_493 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_493;

architecture SYN_BEHAVIORAL of FA_493 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_492 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_492;

architecture SYN_BEHAVIORAL of FA_492 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_491 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_491;

architecture SYN_BEHAVIORAL of FA_491 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_490 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_490;

architecture SYN_BEHAVIORAL of FA_490 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_489 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_489;

architecture SYN_BEHAVIORAL of FA_489 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_488 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_488;

architecture SYN_BEHAVIORAL of FA_488 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_487 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_487;

architecture SYN_BEHAVIORAL of FA_487 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_486 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_486;

architecture SYN_BEHAVIORAL of FA_486 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_485 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_485;

architecture SYN_BEHAVIORAL of FA_485 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_484;

architecture SYN_BEHAVIORAL of FA_484 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_483;

architecture SYN_BEHAVIORAL of FA_483 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_482 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_482;

architecture SYN_BEHAVIORAL of FA_482 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_481;

architecture SYN_BEHAVIORAL of FA_481 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_480 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_480;

architecture SYN_BEHAVIORAL of FA_480 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_479 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_479;

architecture SYN_BEHAVIORAL of FA_479 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_478 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_478;

architecture SYN_BEHAVIORAL of FA_478 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_477 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_477;

architecture SYN_BEHAVIORAL of FA_477 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_476 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_476;

architecture SYN_BEHAVIORAL of FA_476 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_475 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_475;

architecture SYN_BEHAVIORAL of FA_475 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_474 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_474;

architecture SYN_BEHAVIORAL of FA_474 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_473 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_473;

architecture SYN_BEHAVIORAL of FA_473 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_472 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_472;

architecture SYN_BEHAVIORAL of FA_472 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_471 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_471;

architecture SYN_BEHAVIORAL of FA_471 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => Ci, B => A, Z => n3);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_470 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_470;

architecture SYN_BEHAVIORAL of FA_470 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_469 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_469;

architecture SYN_BEHAVIORAL of FA_469 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_468 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_468;

architecture SYN_BEHAVIORAL of FA_468 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => Ci, B => A, Z => n3);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_467 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_467;

architecture SYN_BEHAVIORAL of FA_467 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_466 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_466;

architecture SYN_BEHAVIORAL of FA_466 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_465 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_465;

architecture SYN_BEHAVIORAL of FA_465 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_464;

architecture SYN_BEHAVIORAL of FA_464 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_463;

architecture SYN_BEHAVIORAL of FA_463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => A, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_462;

architecture SYN_BEHAVIORAL of FA_462 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_461;

architecture SYN_BEHAVIORAL of FA_461 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_460;

architecture SYN_BEHAVIORAL of FA_460 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_459;

architecture SYN_BEHAVIORAL of FA_459 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_458;

architecture SYN_BEHAVIORAL of FA_458 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X2 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_457;

architecture SYN_BEHAVIORAL of FA_457 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => A, Z => n1);
   U2 : XOR2_X1 port map( A => n1, B => n2, Z => S);
   U3 : XOR2_X1 port map( A => B, B => Ci, Z => n2);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => Co);
   U7 : NAND2_X1 port map( A1 => n1, A2 => B, ZN => n7);
   U8 : XNOR2_X1 port map( A => n6, B => n5, ZN => n8);
   U9 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U10 : INV_X1 port map( A => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_456;

architecture SYN_BEHAVIORAL of FA_456 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_455;

architecture SYN_BEHAVIORAL of FA_455 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_454;

architecture SYN_BEHAVIORAL of FA_454 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_453;

architecture SYN_BEHAVIORAL of FA_453 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n_1034 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : INV_X1 port map( A => B, ZN => n2);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U5 : FA_X1 port map( A => Ci, B => B, CI => A, CO => n_1034, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_452;

architecture SYN_BEHAVIORAL of FA_452 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_451;

architecture SYN_BEHAVIORAL of FA_451 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NOR2_X2 port map( A1 => n4, A2 => n3, ZN => Co);
   U2 : BUF_X1 port map( A => A, Z => n1);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U5 : AOI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n4);
   U6 : NOR2_X1 port map( A1 => B, A2 => n1, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_450;

architecture SYN_BEHAVIORAL of FA_450 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n1, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n1, B2 => B, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_449;

architecture SYN_BEHAVIORAL of FA_449 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28344, net28345, net28348, net33793, n1, n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : INV_X1 port map( A => B, ZN => net28345);
   U4 : INV_X1 port map( A => A, ZN => net28344);
   U5 : AND2_X1 port map( A1 => net28344, A2 => Ci, ZN => net28348);
   U6 : AND2_X1 port map( A1 => Ci, A2 => net28345, ZN => net33793);
   U7 : XNOR2_X1 port map( A => net33793, B => net28348, ZN => n2);
   U8 : OAI21_X1 port map( B1 => net28344, B2 => net28345, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_448;

architecture SYN_BEHAVIORAL of FA_448 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => B, Z => n1);
   U2 : AOI22_X2 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => n6, B => n1, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U8 : INV_X1 port map( A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_447;

architecture SYN_BEHAVIORAL of FA_447 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28334, net28335, net28336, net28337, net34016, net34415, n1 : 
      std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : CLKBUF_X1 port map( A => A, Z => net34415);
   U4 : CLKBUF_X1 port map( A => Ci, Z => net34016);
   U5 : NAND2_X1 port map( A1 => B, A2 => net34415, ZN => net28334);
   U6 : INV_X1 port map( A => B, ZN => net28337);
   U7 : INV_X1 port map( A => net34016, ZN => net28335);
   U8 : INV_X1 port map( A => net34415, ZN => net28336);
   U9 : AOI22_X1 port map( A1 => net28334, A2 => net28335, B1 => net28336, B2 
                           => net28337, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_446;

architecture SYN_BEHAVIORAL of FA_446 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U3 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_445;

architecture SYN_BEHAVIORAL of FA_445 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28326, net28327, net28328, net28329, n1 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => net28326, A2 => net28327, B1 => net28328, B2 
                           => net28329, ZN => Co);
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net28326);
   U5 : INV_X1 port map( A => B, ZN => net28329);
   U6 : INV_X1 port map( A => Ci, ZN => net28327);
   U7 : INV_X1 port map( A => A, ZN => net28328);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_444;

architecture SYN_BEHAVIORAL of FA_444 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U3 : INV_X1 port map( A => n5, ZN => n2);
   U4 : XNOR2_X1 port map( A => Ci, B => A, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => n2, A => n1, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_443;

architecture SYN_BEHAVIORAL of FA_443 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_442;

architecture SYN_BEHAVIORAL of FA_442 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X2 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U5 : INV_X1 port map( A => Ci, ZN => n2);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_441;

architecture SYN_BEHAVIORAL of FA_441 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_440;

architecture SYN_BEHAVIORAL of FA_440 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_439;

architecture SYN_BEHAVIORAL of FA_439 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_438;

architecture SYN_BEHAVIORAL of FA_438 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n1, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_437;

architecture SYN_BEHAVIORAL of FA_437 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U3 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U4 : INV_X1 port map( A => n1, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_436;

architecture SYN_BEHAVIORAL of FA_436 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n_1035 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : INV_X1 port map( A => B, ZN => n2);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U5 : FA_X1 port map( A => B, B => Ci, CI => A, CO => n_1035, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_435;

architecture SYN_BEHAVIORAL of FA_435 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_434;

architecture SYN_BEHAVIORAL of FA_434 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_433;

architecture SYN_BEHAVIORAL of FA_433 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n3);
   U3 : INV_X1 port map( A => B, ZN => n2);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n4);
   U5 : INV_X1 port map( A => Ci, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n2, B1 => n4, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_432;

architecture SYN_BEHAVIORAL of FA_432 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_431;

architecture SYN_BEHAVIORAL of FA_431 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_430;

architecture SYN_BEHAVIORAL of FA_430 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_429;

architecture SYN_BEHAVIORAL of FA_429 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_428 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_428;

architecture SYN_BEHAVIORAL of FA_428 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_427 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_427;

architecture SYN_BEHAVIORAL of FA_427 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_426 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_426;

architecture SYN_BEHAVIORAL of FA_426 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_425 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_425;

architecture SYN_BEHAVIORAL of FA_425 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_424 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_424;

architecture SYN_BEHAVIORAL of FA_424 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_423 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_423;

architecture SYN_BEHAVIORAL of FA_423 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_422 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_422;

architecture SYN_BEHAVIORAL of FA_422 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_421 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_421;

architecture SYN_BEHAVIORAL of FA_421 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_420;

architecture SYN_BEHAVIORAL of FA_420 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n3, Z => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n1, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_419;

architecture SYN_BEHAVIORAL of FA_419 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_418;

architecture SYN_BEHAVIORAL of FA_418 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_417;

architecture SYN_BEHAVIORAL of FA_417 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_416;

architecture SYN_BEHAVIORAL of FA_416 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_415;

architecture SYN_BEHAVIORAL of FA_415 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_414;

architecture SYN_BEHAVIORAL of FA_414 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_413;

architecture SYN_BEHAVIORAL of FA_413 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_412;

architecture SYN_BEHAVIORAL of FA_412 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => n1, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_411;

architecture SYN_BEHAVIORAL of FA_411 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_410;

architecture SYN_BEHAVIORAL of FA_410 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U3 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => n1, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n1, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_409;

architecture SYN_BEHAVIORAL of FA_409 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_408;

architecture SYN_BEHAVIORAL of FA_408 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_407;

architecture SYN_BEHAVIORAL of FA_407 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_406;

architecture SYN_BEHAVIORAL of FA_406 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_405;

architecture SYN_BEHAVIORAL of FA_405 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_404;

architecture SYN_BEHAVIORAL of FA_404 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_403;

architecture SYN_BEHAVIORAL of FA_403 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_402;

architecture SYN_BEHAVIORAL of FA_402 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : XNOR2_X1 port map( A => A, B => n6, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n6);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => A, ZN => n3);
   U7 : INV_X1 port map( A => n1, ZN => n2);
   U8 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_401;

architecture SYN_BEHAVIORAL of FA_401 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_400;

architecture SYN_BEHAVIORAL of FA_400 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => n1, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n1, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_399;

architecture SYN_BEHAVIORAL of FA_399 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_398;

architecture SYN_BEHAVIORAL of FA_398 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28155, net28156, net28157, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U3 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => net28157);
   U4 : INV_X1 port map( A => B, ZN => net28156);
   U5 : INV_X1 port map( A => A, ZN => net28155);
   U6 : OAI21_X1 port map( B1 => net28155, B2 => net28156, A => net28157, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_397;

architecture SYN_BEHAVIORAL of FA_397 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => Ci, B => B, Z => n3);
   U5 : XOR2_X1 port map( A => A, B => n3, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_396;

architecture SYN_BEHAVIORAL of FA_396 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_395;

architecture SYN_BEHAVIORAL of FA_395 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_394;

architecture SYN_BEHAVIORAL of FA_394 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_393;

architecture SYN_BEHAVIORAL of FA_393 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_392;

architecture SYN_BEHAVIORAL of FA_392 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_391;

architecture SYN_BEHAVIORAL of FA_391 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_390 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_390;

architecture SYN_BEHAVIORAL of FA_390 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_389 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_389;

architecture SYN_BEHAVIORAL of FA_389 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_388 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_388;

architecture SYN_BEHAVIORAL of FA_388 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_387;

architecture SYN_BEHAVIORAL of FA_387 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_386 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_386;

architecture SYN_BEHAVIORAL of FA_386 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_385 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_385;

architecture SYN_BEHAVIORAL of FA_385 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_384 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_384;

architecture SYN_BEHAVIORAL of FA_384 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_383 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_383;

architecture SYN_BEHAVIORAL of FA_383 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_382 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_382;

architecture SYN_BEHAVIORAL of FA_382 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_381 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_381;

architecture SYN_BEHAVIORAL of FA_381 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_380;

architecture SYN_BEHAVIORAL of FA_380 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_379;

architecture SYN_BEHAVIORAL of FA_379 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_378 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_378;

architecture SYN_BEHAVIORAL of FA_378 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_377;

architecture SYN_BEHAVIORAL of FA_377 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_376;

architecture SYN_BEHAVIORAL of FA_376 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_375;

architecture SYN_BEHAVIORAL of FA_375 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_374;

architecture SYN_BEHAVIORAL of FA_374 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_373;

architecture SYN_BEHAVIORAL of FA_373 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_372;

architecture SYN_BEHAVIORAL of FA_372 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_371;

architecture SYN_BEHAVIORAL of FA_371 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_370;

architecture SYN_BEHAVIORAL of FA_370 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_369;

architecture SYN_BEHAVIORAL of FA_369 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_368;

architecture SYN_BEHAVIORAL of FA_368 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => B, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_367;

architecture SYN_BEHAVIORAL of FA_367 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_366;

architecture SYN_BEHAVIORAL of FA_366 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_365 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_365;

architecture SYN_BEHAVIORAL of FA_365 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_364 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_364;

architecture SYN_BEHAVIORAL of FA_364 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_363 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_363;

architecture SYN_BEHAVIORAL of FA_363 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_362 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_362;

architecture SYN_BEHAVIORAL of FA_362 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_361 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_361;

architecture SYN_BEHAVIORAL of FA_361 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_360 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_360;

architecture SYN_BEHAVIORAL of FA_360 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_359 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_359;

architecture SYN_BEHAVIORAL of FA_359 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_358 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_358;

architecture SYN_BEHAVIORAL of FA_358 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_357 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_357;

architecture SYN_BEHAVIORAL of FA_357 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_356 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_356;

architecture SYN_BEHAVIORAL of FA_356 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : INV_X1 port map( A => B, ZN => n2);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U5 : XOR2_X1 port map( A => Ci, B => B, Z => n4);
   U6 : XOR2_X1 port map( A => A, B => n4, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_355 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_355;

architecture SYN_BEHAVIORAL of FA_355 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_354 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_354;

architecture SYN_BEHAVIORAL of FA_354 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_353 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_353;

architecture SYN_BEHAVIORAL of FA_353 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_352 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_352;

architecture SYN_BEHAVIORAL of FA_352 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_351 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_351;

architecture SYN_BEHAVIORAL of FA_351 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_350 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_350;

architecture SYN_BEHAVIORAL of FA_350 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_349 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_349;

architecture SYN_BEHAVIORAL of FA_349 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_348 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_348;

architecture SYN_BEHAVIORAL of FA_348 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_347 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_347;

architecture SYN_BEHAVIORAL of FA_347 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_346 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_346;

architecture SYN_BEHAVIORAL of FA_346 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_345 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_345;

architecture SYN_BEHAVIORAL of FA_345 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_344;

architecture SYN_BEHAVIORAL of FA_344 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_343;

architecture SYN_BEHAVIORAL of FA_343 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_342;

architecture SYN_BEHAVIORAL of FA_342 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_341;

architecture SYN_BEHAVIORAL of FA_341 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_340;

architecture SYN_BEHAVIORAL of FA_340 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_339;

architecture SYN_BEHAVIORAL of FA_339 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U5 : XOR2_X1 port map( A => Ci, B => B, Z => n4);
   U6 : XOR2_X1 port map( A => n1, B => n4, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_338;

architecture SYN_BEHAVIORAL of FA_338 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_337;

architecture SYN_BEHAVIORAL of FA_337 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_336;

architecture SYN_BEHAVIORAL of FA_336 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => B, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_335;

architecture SYN_BEHAVIORAL of FA_335 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_334;

architecture SYN_BEHAVIORAL of FA_334 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => B, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_333;

architecture SYN_BEHAVIORAL of FA_333 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_332;

architecture SYN_BEHAVIORAL of FA_332 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_331;

architecture SYN_BEHAVIORAL of FA_331 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_330;

architecture SYN_BEHAVIORAL of FA_330 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n_1036 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => A, Z => n1);
   U2 : INV_X1 port map( A => n1, ZN => n4);
   U3 : INV_X1 port map( A => B, ZN => n3);
   U4 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U6 : FA_X1 port map( A => Ci, B => B, CI => A, CO => n_1036, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_329;

architecture SYN_BEHAVIORAL of FA_329 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_328;

architecture SYN_BEHAVIORAL of FA_328 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n2);
   U2 : CLKBUF_X1 port map( A => A, Z => n1);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n6);
   U4 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : INV_X1 port map( A => n1, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n1, B2 => B, A => n2, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_327;

architecture SYN_BEHAVIORAL of FA_327 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_326;

architecture SYN_BEHAVIORAL of FA_326 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => A, Z => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U5 : XOR2_X1 port map( A => Ci, B => B, Z => n4);
   U6 : XOR2_X1 port map( A => n1, B => n4, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_325;

architecture SYN_BEHAVIORAL of FA_325 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27876, net27877, net27878, net27879, net34482, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net27878);
   U4 : INV_X1 port map( A => B, ZN => net27877);
   U5 : CLKBUF_X1 port map( A => A, Z => net34482);
   U6 : INV_X1 port map( A => Ci, ZN => net27879);
   U7 : AOI22_X2 port map( A1 => net27876, A2 => net27877, B1 => net27878, B2 
                           => net27879, ZN => Co);
   U8 : INV_X1 port map( A => net34482, ZN => net27876);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_324;

architecture SYN_BEHAVIORAL of FA_324 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n1);
   U2 : NAND2_X1 port map( A1 => n1, A2 => n7, ZN => n2);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n3);
   U4 : AND2_X2 port map( A1 => n3, A2 => n2, ZN => Co);
   U5 : INV_X1 port map( A => n8, ZN => n4);
   U6 : XNOR2_X1 port map( A => A, B => Ci, ZN => n9);
   U7 : XNOR2_X1 port map( A => n9, B => B, ZN => S);
   U8 : INV_X1 port map( A => A, ZN => n8);
   U9 : INV_X1 port map( A => B, ZN => n7);
   U10 : NAND2_X1 port map( A1 => B, A2 => n4, ZN => n6);
   U11 : INV_X1 port map( A => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_323;

architecture SYN_BEHAVIORAL of FA_323 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net35527, net35526, net35530, n1 : std_logic;

begin
   
   U1 : NOR2_X2 port map( A1 => net35527, A2 => net35526, ZN => Co);
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U4 : BUF_X1 port map( A => A, Z => net35530);
   U5 : AOI21_X1 port map( B1 => net35530, B2 => Ci, A => B, ZN => net35527);
   U6 : NOR2_X1 port map( A1 => net35530, A2 => Ci, ZN => net35526);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_322;

architecture SYN_BEHAVIORAL of FA_322 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : AOI22_X2 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U3 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U7 : INV_X1 port map( A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_321;

architecture SYN_BEHAVIORAL of FA_321 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27856, net27857, net27858, net27859, net34519, n1, n2 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => net27856, A2 => net27857, B1 => net27858, B2 
                           => net27859, ZN => Co);
   U2 : CLKBUF_X1 port map( A => B, Z => n1);
   U3 : INV_X1 port map( A => A, ZN => net27858);
   U4 : XNOR2_X1 port map( A => Ci, B => B, ZN => n2);
   U5 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => net27856);
   U6 : INV_X1 port map( A => n1, ZN => net27859);
   U7 : XNOR2_X1 port map( A => n2, B => A, ZN => S);
   U8 : CLKBUF_X1 port map( A => Ci, Z => net34519);
   U9 : INV_X1 port map( A => net34519, ZN => net27857);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_320;

architecture SYN_BEHAVIORAL of FA_320 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);
   U2 : BUF_X1 port map( A => B, Z => n1);
   U3 : XNOR2_X1 port map( A => n2, B => n1, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => A, ZN => n4);
   U8 : INV_X1 port map( A => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_319;

architecture SYN_BEHAVIORAL of FA_319 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_318;

architecture SYN_BEHAVIORAL of FA_318 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : AOI22_X2 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U3 : XNOR2_X1 port map( A => n6, B => A, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U6 : INV_X1 port map( A => n1, ZN => n4);
   U7 : INV_X1 port map( A => A, ZN => n3);
   U8 : INV_X1 port map( A => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_317;

architecture SYN_BEHAVIORAL of FA_317 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n1);
   U2 : AOI21_X2 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => n5, B => n1, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net27835, net27836, net27837, n1, n2 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n2);
   U3 : XNOR2_X1 port map( A => A, B => n2, ZN => S);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => n1, ZN => net27837);
   U5 : INV_X1 port map( A => B, ZN => net27836);
   U6 : INV_X1 port map( A => A, ZN => net27835);
   U7 : OAI21_X1 port map( B1 => net27835, B2 => net27836, A => net27837, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => n1, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => Ci, B => A, Z => n3);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_304;

architecture SYN_BEHAVIORAL of FA_304 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_303;

architecture SYN_BEHAVIORAL of FA_303 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_302;

architecture SYN_BEHAVIORAL of FA_302 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_301;

architecture SYN_BEHAVIORAL of FA_301 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_300;

architecture SYN_BEHAVIORAL of FA_300 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_299;

architecture SYN_BEHAVIORAL of FA_299 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_298;

architecture SYN_BEHAVIORAL of FA_298 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_297;

architecture SYN_BEHAVIORAL of FA_297 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_296;

architecture SYN_BEHAVIORAL of FA_296 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_295;

architecture SYN_BEHAVIORAL of FA_295 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_294;

architecture SYN_BEHAVIORAL of FA_294 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_293;

architecture SYN_BEHAVIORAL of FA_293 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : CLKBUF_X1 port map( A => n6, Z => n2);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U4 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => n1, ZN => n3);
   U8 : OAI22_X1 port map( A1 => n2, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n1);
   U2 : INV_X1 port map( A => n5, ZN => n2);
   U3 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => n2, A => n1, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : INV_X1 port map( A => n5, ZN => n2);
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n1, B2 => n2, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X4
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI222_X4 port map( A1 => n3, A2 => n2, B1 => n1, B2 => n2, C1 => n1, 
                           C2 => n3, ZN => Co);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net27515, net31517, net34434, n1, n2 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => A, Z => net31517);
   U2 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U4 : OAI21_X1 port map( B1 => net31517, B2 => net34434, A => Ci, ZN => 
                           net27515);
   U5 : CLKBUF_X1 port map( A => B, Z => net34434);
   U6 : NAND2_X1 port map( A1 => net27515, A2 => n2, ZN => Co);
   U7 : NAND2_X1 port map( A1 => net31517, A2 => net34434, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => A, Z => n1);
   U2 : AOI22_X2 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U5 : INV_X1 port map( A => n1, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : NAND2_X1 port map( A1 => B, A2 => n1, ZN => n3);
   U8 : INV_X1 port map( A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27506, net27507, net27508, net34815, net42254, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : CLKBUF_X1 port map( A => Ci, Z => net42254);
   U4 : INV_X1 port map( A => A, ZN => net27506);
   U5 : OAI21_X1 port map( B1 => B, B2 => net34815, A => net42254, ZN => 
                           net27508);
   U6 : INV_X1 port map( A => B, ZN => net27507);
   U7 : INV_X1 port map( A => net27506, ZN => net34815);
   U8 : OAI21_X1 port map( B1 => net27506, B2 => net27507, A => net27508, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27501, net27502, net27503, net27504, net34834, n1, n2, n3 : 
      std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => A, A2 => net34834, ZN => net27503);
   U4 : INV_X1 port map( A => A, ZN => net27501);
   U5 : INV_X1 port map( A => B, ZN => net27502);
   U6 : INV_X1 port map( A => Ci, ZN => net27504);
   U7 : NAND2_X1 port map( A1 => net27501, A2 => net27502, ZN => n2);
   U8 : NAND2_X1 port map( A1 => net27503, A2 => net27504, ZN => n3);
   U9 : AND2_X2 port map( A1 => n2, A2 => n3, ZN => Co);
   U10 : INV_X1 port map( A => net27502, ZN => net34834);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net27497, net27498, net27499, n1, n2 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => net27498);
   U5 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => net27499);
   U6 : INV_X1 port map( A => n1, ZN => net27497);
   U7 : OAI21_X1 port map( B1 => net27497, B2 => net27498, A => net27499, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n_1037 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n2);
   U3 : AND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);
   U4 : CLKBUF_X1 port map( A => B, Z => n3);
   U5 : INV_X1 port map( A => n6, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => n8);
   U7 : INV_X1 port map( A => Ci, ZN => n7);
   U8 : INV_X1 port map( A => A, ZN => n6);
   U9 : INV_X1 port map( A => n3, ZN => n5);
   U10 : FA_X1 port map( A => B, B => Ci, CI => A, CO => n_1037, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => n1);
   U2 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n1, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U6 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X2 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27478, net27476, n1, n2 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n1, B2 => net27478, A => n2, ZN => Co);
   U2 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => net27476);
   U5 : INV_X1 port map( A => Ci, ZN => net27478);
   U6 : XNOR2_X1 port map( A => Ci, B => net27476, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X2 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : INV_X1 port map( A => Ci, ZN => n2);
   U3 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U5 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U6 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n_1038 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : INV_X1 port map( A => B, ZN => n2);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U5 : FA_X1 port map( A => Ci, B => A, CI => B, CO => n_1038, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n2);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n2, ZN => S);
   U5 : INV_X1 port map( A => n1, ZN => n4);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => B, ZN => n3);
   U8 : OAI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n1);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n1, ZN => n3);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => n1, Z => S);
   U2 : XOR2_X1 port map( A => Ci, B => A, Z => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X2 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => n3, A2 => n4, ZN => n1);
   U2 : NAND2_X2 port map( A1 => n1, A2 => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n3);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U3 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U4 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n3);
   U7 : OAI21_X1 port map( B1 => n1, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27323, net27324, net27325, n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => net27323, ZN => n1);
   U2 : OAI21_X2 port map( B1 => net27323, B2 => net27324, A => net27325, ZN =>
                           Co);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => net27324);
   U6 : OAI21_X1 port map( B1 => n1, B2 => B, A => Ci, ZN => net27325);
   U7 : INV_X1 port map( A => A, ZN => net27323);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => n2, B => A, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => Ci, ZN => n2);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => n1, ZN => n4);
   U7 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27315, net27316, net27317, net31457, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : BUF_X1 port map( A => A, Z => net31457);
   U4 : OAI21_X1 port map( B1 => net31457, B2 => B, A => Ci, ZN => net27317);
   U5 : INV_X1 port map( A => B, ZN => net27316);
   U6 : OAI21_X1 port map( B1 => net27315, B2 => net27316, A => net27317, ZN =>
                           Co);
   U7 : INV_X1 port map( A => net31457, ZN => net27315);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net27312, net27313, n1, n2, n3 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n1);
   U3 : XNOR2_X1 port map( A => n2, B => n1, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net27312);
   U6 : NAND2_X1 port map( A1 => n3, A2 => B, ZN => net27313);
   U7 : NAND2_X1 port map( A1 => net27313, A2 => net27312, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27308, net27309, net27310, net34232, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : INV_X1 port map( A => B, ZN => net27309);
   U4 : CLKBUF_X1 port map( A => A, Z => net34232);
   U5 : OAI21_X1 port map( B1 => B, B2 => net34232, A => Ci, ZN => net27310);
   U6 : INV_X1 port map( A => net34232, ZN => net27308);
   U7 : OAI21_X1 port map( B1 => net27308, B2 => net27309, A => net27310, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n3);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => Co);
   U3 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U5 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => B, ZN => n2);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => Co);
   U3 : INV_X1 port map( A => n4, ZN => n1);
   U4 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U6 : INV_X1 port map( A => A, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n1);
   U2 : XNOR2_X1 port map( A => n4, B => n1, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : OAI21_X2 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   U2 : CLKBUF_X1 port map( A => B, Z => n1);
   U3 : INV_X1 port map( A => n5, ZN => n2);
   U4 : XNOR2_X1 port map( A => A, B => n6, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => Ci, ZN => n6);
   U6 : INV_X1 port map( A => A, ZN => n5);
   U7 : INV_X1 port map( A => n1, ZN => n4);
   U8 : OAI21_X1 port map( B1 => n1, B2 => n2, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27284, net27285, net27286, n1, n2, n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => net27284, ZN => n1);
   U2 : OAI21_X1 port map( B1 => net27284, B2 => net27285, A => net27286, ZN =>
                           Co);
   U3 : INV_X1 port map( A => net27285, ZN => n2);
   U4 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U5 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U6 : OAI21_X1 port map( B1 => n2, B2 => n1, A => Ci, ZN => net27286);
   U7 : INV_X1 port map( A => B, ZN => net27285);
   U8 : INV_X1 port map( A => A, ZN => net27284);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => B, Z => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => n4, B => n1, ZN => S);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U6 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => n1);
   U2 : INV_X1 port map( A => n4, ZN => n2);
   U3 : XNOR2_X1 port map( A => n6, B => A, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => B, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => n2, B2 => n1, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI22_X2 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => n1);
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL_architecture of FA_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL_architecture2 of FA_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL_architecture3 of FA_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL_architecture of FA_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL_architecture2 of FA_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL_architecture3 of FA_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL_architecture of FA_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL_architecture2 of FA_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL_architecture3 of FA_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL_architecture of FA_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL_architecture2 of FA_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL_architecture3 of FA_109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL_architecture of FA_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL_architecture2 of FA_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL_architecture3 of FA_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL_architecture of FA_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL_architecture2 of FA_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL_architecture3 of FA_101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL_architecture of FA_99 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL_architecture2 of FA_98 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL_architecture3 of FA_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL_architecture of FA_95 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL_architecture2 of FA_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL_architecture3 of FA_93 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL_architecture of FA_91 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL_architecture2 of FA_90 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL_architecture3 of FA_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL_architecture of FA_87 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL_architecture2 of FA_86 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL_architecture3 of FA_85 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n3, Z => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n1, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL_architecture of FA_83 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL_architecture2 of FA_82 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL_architecture3 of FA_81 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => n1, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL_architecture of FA_79 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL_architecture2 of FA_78 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL_architecture3 of FA_77 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n3, Z => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n1, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL_architecture of FA_75 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n1);
   U2 : INV_X1 port map( A => A, ZN => n3);
   U3 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n3, B2 => n2, ZN => Co);
   U7 : INV_X1 port map( A => n5, ZN => n6);
   U8 : XOR2_X1 port map( A => n1, B => n6, Z => S);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL_architecture2 of FA_74 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL_architecture3 of FA_73 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => n1, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL_architecture of FA_71 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL_architecture2 of FA_70 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL_architecture3 of FA_69 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n3, Z => n1);
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n1, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL_architecture of FA_67 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL_architecture2 of FA_66 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL_architecture3 of FA_65 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n1);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => n1, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL_architecture of FA_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL_architecture2 of FA_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL_architecture3 of FA_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => Ci, B => A, Z => n3);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL_architecture of FA_59 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL_architecture2 of FA_58 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL_architecture3 of FA_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL_architecture of FA_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL_architecture2 of FA_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL_architecture3 of FA_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : XOR2_X1 port map( A => Ci, B => A, Z => n3);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL_architecture of FA_51 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL_architecture2 of FA_50 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL_architecture3 of FA_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL_architecture of FA_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL_architecture2 of FA_46 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL_architecture3 of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : INV_X1 port map( A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U5 : XOR2_X1 port map( A => A, B => Ci, Z => n4);
   U6 : XOR2_X1 port map( A => B, B => n4, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL_architecture of FA_43 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL_architecture2 of FA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL_architecture3 of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL_architecture of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL_architecture2 of FA_38 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL_architecture3 of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : XOR2_X1 port map( A => Ci, B => A, Z => n3);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL_architecture of FA_35 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL_architecture2 of FA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL_architecture3 of FA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL_architecture of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL_architecture2 of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL_architecture3 of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL_architecture of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL_architecture2 of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL_architecture3 of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL_architecture of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL_architecture2 of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL_architecture3 of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL_architecture of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL_architecture2 of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL_architecture3 of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL_architecture of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL_architecture2 of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL_architecture3 of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL_architecture of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL_architecture2 of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL_architecture3 of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL_architecture of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL_architecture2 of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL_architecture3 of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL_architecture of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL_architecture2 of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL_architecture3 of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_43 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_43;

architecture SYN_rtl of HA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X2 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_42 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_42;

architecture SYN_rtl of HA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_41 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_41;

architecture SYN_rtl of HA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_40 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_40;

architecture SYN_rtl of HA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_39 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_39;

architecture SYN_rtl of HA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_38 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_38;

architecture SYN_rtl of HA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_37 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_37;

architecture SYN_rtl of HA_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => n2, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => S);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_36 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_36;

architecture SYN_rtl of HA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_35 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_35;

architecture SYN_rtl of HA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_34 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_34;

architecture SYN_rtl of HA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_33 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_33;

architecture SYN_rtl of HA_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => S);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : INV_X1 port map( A => A, ZN => n2);
   U5 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U6 : NAND2_X1 port map( A1 => B, A2 => n2, ZN => n3);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_32 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_32;

architecture SYN_rtl of HA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_31 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_31;

architecture SYN_rtl of HA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_30 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_30;

architecture SYN_rtl of HA_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_29 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_29;

architecture SYN_rtl of HA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_28 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_28;

architecture SYN_rtl of HA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_27 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_27;

architecture SYN_rtl of HA_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_26 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_26;

architecture SYN_rtl of HA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_25 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_25;

architecture SYN_rtl of HA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_24 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_24;

architecture SYN_rtl of HA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_23 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_23;

architecture SYN_rtl of HA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_22 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_22;

architecture SYN_rtl of HA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_21 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_21;

architecture SYN_rtl of HA_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : INV_X1 port map( A => B, ZN => n1);
   U3 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => C);
   U4 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_20 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_20;

architecture SYN_rtl of HA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_19 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_19;

architecture SYN_rtl of HA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_18 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_18;

architecture SYN_rtl of HA_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_17 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_17;

architecture SYN_rtl of HA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_16 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_16;

architecture SYN_rtl of HA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_15 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_15;

architecture SYN_rtl of HA_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_14 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_14;

architecture SYN_rtl of HA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_13 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_13;

architecture SYN_rtl of HA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_12 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_12;

architecture SYN_rtl of HA_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_11 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_11;

architecture SYN_rtl of HA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_10 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_10;

architecture SYN_rtl of HA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_9 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_9;

architecture SYN_rtl of HA_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_8 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_8;

architecture SYN_rtl of HA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_7 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_7;

architecture SYN_rtl of HA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_6 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_6;

architecture SYN_rtl of HA_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_5 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_5;

architecture SYN_rtl of HA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_4 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_4;

architecture SYN_rtl of HA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_3 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_3;

architecture SYN_rtl of HA_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_2 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_2;

architecture SYN_rtl of HA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_1 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_1;

architecture SYN_rtl of HA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_16 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_16;

architecture SYN_beh of ENC_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A(27), ZN => n4);
   U4 : CLKBUF_X1 port map( A => b(1), Z => n1);
   U5 : CLKBUF_X1 port map( A => b(2), Z => n2);
   U6 : CLKBUF_X1 port map( A => b(2), Z => n15);
   U7 : BUF_X1 port map( A => b(0), Z => n6);
   U8 : BUF_X1 port map( A => n102, Z => n24);
   U9 : CLKBUF_X1 port map( A => n102, Z => n8);
   U10 : BUF_X2 port map( A => n100, Z => n16);
   U11 : NAND2_X1 port map( A1 => n12, A2 => n2, ZN => n3);
   U12 : MUX2_X1 port map( A => n98, B => n3, S => n4, Z => n88);
   U13 : NAND2_X1 port map( A1 => n62, A2 => n2, ZN => n5);
   U14 : NAND2_X1 port map( A1 => n62, A2 => n2, ZN => n104);
   U15 : CLKBUF_X1 port map( A => n104, Z => n26);
   U16 : BUF_X1 port map( A => n100, Z => n18);
   U17 : INV_X1 port map( A => b(0), ZN => n7);
   U18 : BUF_X2 port map( A => n5, Z => n25);
   U19 : INV_X1 port map( A => b(1), ZN => n9);
   U20 : BUF_X1 port map( A => n102, Z => n22);
   U21 : NAND2_X1 port map( A1 => n6, A2 => n1, ZN => n10);
   U22 : BUF_X2 port map( A => n10, Z => n19);
   U23 : BUF_X2 port map( A => n100, Z => n17);
   U24 : CLKBUF_X1 port map( A => n10, Z => n21);
   U25 : BUF_X1 port map( A => n102, Z => n23);
   U26 : BUF_X1 port map( A => n10, Z => n20);
   U27 : XNOR2_X1 port map( A => b(0), B => n9, ZN => n11);
   U28 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => n12);
   U29 : NAND2_X1 port map( A1 => n11, A2 => n63, ZN => n13);
   U30 : NAND2_X1 port map( A1 => n11, A2 => n63, ZN => n95);
   U31 : NAND2_X1 port map( A1 => n11, A2 => n63, ZN => n69);
   U32 : CLKBUF_X1 port map( A => n5, Z => n14);
   U33 : INV_X1 port map( A => n15, ZN => n63);
   U34 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n28);
   U35 : INV_X1 port map( A => b(1), ZN => n31);
   U36 : INV_X1 port map( A => b(0), ZN => n30);
   U37 : NAND3_X1 port map( A1 => n7, A2 => n31, A3 => b(2), ZN => n102);
   U38 : NAND2_X1 port map( A1 => n28, A2 => b(2), ZN => n29);
   U39 : MUX2_X1 port map( A => n29, B => n13, S => A(0), Z => n27);
   U40 : OAI211_X1 port map( C1 => n63, C2 => n10, A => n23, B => n27, ZN => 
                           p(0));
   U41 : MUX2_X1 port map( A => n8, B => n21, S => A(0), Z => n33);
   U42 : NAND2_X1 port map( A1 => n29, A2 => n15, ZN => n100);
   U43 : NAND2_X1 port map( A1 => n30, A2 => n9, ZN => n62);
   U44 : MUX2_X1 port map( A => n25, B => n13, S => A(1), Z => n32);
   U45 : NAND3_X1 port map( A1 => n33, A2 => n17, A3 => n32, ZN => p(1));
   U46 : MUX2_X1 port map( A => n8, B => n21, S => A(1), Z => n35);
   U47 : MUX2_X1 port map( A => n25, B => n13, S => A(2), Z => n34);
   U48 : NAND3_X1 port map( A1 => n35, A2 => n16, A3 => n34, ZN => p(2));
   U49 : MUX2_X1 port map( A => n24, B => n21, S => A(2), Z => n37);
   U50 : MUX2_X1 port map( A => n25, B => n69, S => A(3), Z => n36);
   U51 : NAND3_X1 port map( A1 => n37, A2 => n18, A3 => n36, ZN => p(3));
   U52 : MUX2_X1 port map( A => n23, B => n21, S => A(3), Z => n39);
   U53 : MUX2_X1 port map( A => n25, B => n13, S => A(4), Z => n38);
   U54 : NAND3_X1 port map( A1 => n39, A2 => n17, A3 => n38, ZN => p(4));
   U55 : MUX2_X1 port map( A => n24, B => n21, S => A(4), Z => n41);
   U56 : MUX2_X1 port map( A => n25, B => n69, S => A(5), Z => n40);
   U57 : NAND3_X1 port map( A1 => n41, A2 => n16, A3 => n40, ZN => p(5));
   U58 : MUX2_X1 port map( A => n8, B => n21, S => A(5), Z => n43);
   U59 : MUX2_X1 port map( A => n25, B => n13, S => A(6), Z => n42);
   U60 : NAND3_X1 port map( A1 => n43, A2 => n18, A3 => n42, ZN => p(6));
   U61 : MUX2_X1 port map( A => n24, B => n21, S => A(6), Z => n45);
   U62 : MUX2_X1 port map( A => n25, B => n69, S => A(7), Z => n44);
   U63 : NAND3_X1 port map( A1 => n45, A2 => n17, A3 => n44, ZN => p(7));
   U64 : MUX2_X1 port map( A => n23, B => n21, S => A(7), Z => n47);
   U65 : MUX2_X1 port map( A => n26, B => n13, S => A(8), Z => n46);
   U66 : NAND3_X1 port map( A1 => n47, A2 => n17, A3 => n46, ZN => p(8));
   U67 : MUX2_X1 port map( A => n23, B => n21, S => A(8), Z => n49);
   U68 : MUX2_X1 port map( A => n26, B => n69, S => A(9), Z => n48);
   U69 : NAND3_X1 port map( A1 => n49, A2 => n17, A3 => n48, ZN => p(9));
   U70 : MUX2_X1 port map( A => n24, B => n21, S => A(9), Z => n51);
   U71 : MUX2_X1 port map( A => n5, B => n69, S => A(10), Z => n50);
   U72 : NAND3_X1 port map( A1 => n51, A2 => n18, A3 => n50, ZN => p(10));
   U73 : MUX2_X1 port map( A => n25, B => n13, S => A(11), Z => n53);
   U74 : MUX2_X1 port map( A => n23, B => n20, S => A(10), Z => n52);
   U75 : NAND3_X1 port map( A1 => n53, A2 => n16, A3 => n52, ZN => p(11));
   U76 : MUX2_X1 port map( A => n8, B => n20, S => A(11), Z => n55);
   U77 : MUX2_X1 port map( A => n26, B => n95, S => A(12), Z => n54);
   U78 : NAND3_X1 port map( A1 => n55, A2 => n16, A3 => n54, ZN => p(12));
   U79 : MUX2_X1 port map( A => n14, B => n13, S => A(13), Z => n57);
   U80 : MUX2_X1 port map( A => n24, B => n20, S => A(12), Z => n56);
   U81 : NAND3_X1 port map( A1 => n16, A2 => n57, A3 => n56, ZN => p(13));
   U82 : MUX2_X1 port map( A => n24, B => n20, S => A(13), Z => n59);
   U83 : MUX2_X1 port map( A => n25, B => n13, S => A(14), Z => n58);
   U84 : NAND3_X1 port map( A1 => n59, A2 => n18, A3 => n58, ZN => p(14));
   U85 : MUX2_X1 port map( A => n25, B => n69, S => A(15), Z => n61);
   U86 : MUX2_X1 port map( A => n24, B => n20, S => A(14), Z => n60);
   U87 : NAND3_X1 port map( A1 => n61, A2 => n17, A3 => n60, ZN => p(15));
   U88 : NAND2_X1 port map( A1 => n12, A2 => n15, ZN => n90);
   U89 : XOR2_X1 port map( A => n6, B => n1, Z => n64);
   U90 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => n98);
   U91 : MUX2_X1 port map( A => n25, B => n98, S => A(16), Z => n66);
   U92 : MUX2_X1 port map( A => n23, B => n20, S => A(15), Z => n65);
   U93 : NAND3_X1 port map( A1 => n66, A2 => n17, A3 => n65, ZN => p(16));
   U94 : MUX2_X1 port map( A => n25, B => n98, S => A(17), Z => n68);
   U95 : MUX2_X1 port map( A => n24, B => n20, S => A(16), Z => n67);
   U96 : NAND3_X1 port map( A1 => n68, A2 => n18, A3 => n67, ZN => p(17));
   U97 : MUX2_X1 port map( A => n8, B => n20, S => A(17), Z => n71);
   U98 : MUX2_X1 port map( A => n25, B => n13, S => A(18), Z => n70);
   U99 : NAND3_X1 port map( A1 => n71, A2 => n16, A3 => n70, ZN => p(18));
   U100 : MUX2_X1 port map( A => n3, B => n98, S => A(19), Z => n73);
   U101 : MUX2_X1 port map( A => n24, B => n20, S => A(18), Z => n72);
   U102 : NAND3_X1 port map( A1 => n73, A2 => n16, A3 => n72, ZN => p(19));
   U103 : MUX2_X1 port map( A => n24, B => n20, S => A(19), Z => n75);
   U104 : MUX2_X1 port map( A => n26, B => n69, S => A(20), Z => n74);
   U105 : NAND3_X1 port map( A1 => n75, A2 => n18, A3 => n74, ZN => p(20));
   U106 : MUX2_X1 port map( A => n23, B => n20, S => A(20), Z => n77);
   U107 : MUX2_X1 port map( A => n5, B => n95, S => A(21), Z => n76);
   U108 : NAND3_X1 port map( A1 => n77, A2 => n18, A3 => n76, ZN => p(21));
   U109 : MUX2_X1 port map( A => n24, B => n19, S => A(21), Z => n79);
   U110 : MUX2_X1 port map( A => n90, B => n95, S => A(22), Z => n78);
   U111 : NAND3_X1 port map( A1 => n79, A2 => n16, A3 => n78, ZN => p(22));
   U112 : MUX2_X1 port map( A => n8, B => n19, S => A(22), Z => n81);
   U113 : MUX2_X1 port map( A => n3, B => n95, S => A(23), Z => n80);
   U114 : NAND3_X1 port map( A1 => n81, A2 => n16, A3 => n80, ZN => p(23));
   U115 : MUX2_X1 port map( A => n24, B => n19, S => A(23), Z => n83);
   U116 : MUX2_X1 port map( A => n5, B => n98, S => A(24), Z => n82);
   U117 : NAND3_X1 port map( A1 => n83, A2 => n82, A3 => n18, ZN => p(24));
   U118 : MUX2_X1 port map( A => n22, B => n19, S => A(24), Z => n85);
   U119 : MUX2_X1 port map( A => n90, B => n98, S => A(25), Z => n84);
   U120 : NAND3_X1 port map( A1 => n84, A2 => n85, A3 => n16, ZN => p(25));
   U121 : MUX2_X1 port map( A => n23, B => n19, S => A(25), Z => n87);
   U122 : MUX2_X1 port map( A => n104, B => n98, S => A(26), Z => n86);
   U123 : NAND3_X1 port map( A1 => n87, A2 => n86, A3 => n17, ZN => p(26));
   U124 : MUX2_X1 port map( A => n22, B => n19, S => A(26), Z => n89);
   U125 : NAND3_X1 port map( A1 => n88, A2 => n89, A3 => n17, ZN => p(27));
   U126 : MUX2_X1 port map( A => n22, B => n19, S => A(27), Z => n92);
   U127 : MUX2_X1 port map( A => n90, B => n69, S => A(28), Z => n91);
   U128 : NAND3_X1 port map( A1 => n92, A2 => n17, A3 => n91, ZN => p(28));
   U129 : MUX2_X1 port map( A => n22, B => n19, S => A(28), Z => n94);
   U130 : MUX2_X1 port map( A => n104, B => n69, S => A(29), Z => n93);
   U131 : NAND3_X1 port map( A1 => n93, A2 => n18, A3 => n94, ZN => p(29));
   U132 : MUX2_X1 port map( A => n8, B => n19, S => A(29), Z => n97);
   U133 : MUX2_X1 port map( A => n14, B => n69, S => A(30), Z => n96);
   U134 : NAND3_X1 port map( A1 => n97, A2 => n17, A3 => n96, ZN => p(30));
   U135 : MUX2_X1 port map( A => n8, B => n19, S => A(30), Z => n101);
   U136 : MUX2_X1 port map( A => n25, B => n98, S => A(31), Z => n99);
   U137 : NAND3_X1 port map( A1 => n101, A2 => n18, A3 => n99, ZN => p(31));
   U138 : MUX2_X1 port map( A => n24, B => n19, S => A(31), Z => n103);
   U139 : NAND2_X1 port map( A1 => n25, A2 => n103, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_15 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_15;

architecture SYN_beh of ENC_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101 : 
      std_logic;

begin
   
   U3 : BUF_X1 port map( A => n94, Z => n13);
   U4 : NAND2_X1 port map( A1 => n21, A2 => n61, ZN => n1);
   U5 : INV_X1 port map( A => n61, ZN => n2);
   U6 : AND3_X1 port map( A1 => b(2), A2 => b(0), A3 => b(1), ZN => n3);
   U7 : INV_X1 port map( A => n3, ZN => n96);
   U8 : AND2_X2 port map( A1 => n24, A2 => b(2), ZN => n11);
   U9 : NAND2_X1 port map( A1 => n84, A2 => n4, ZN => n5);
   U10 : NAND2_X1 port map( A1 => n83, A2 => A(23), ZN => n6);
   U11 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => n72);
   U12 : INV_X1 port map( A => A(23), ZN => n4);
   U13 : CLKBUF_X1 port map( A => n14, Z => n7);
   U14 : BUF_X1 port map( A => b(0), Z => n10);
   U15 : NAND2_X1 port map( A1 => n11, A2 => n78, ZN => n93);
   U16 : BUF_X4 port map( A => n101, Z => n20);
   U17 : CLKBUF_X3 port map( A => n96, Z => n15);
   U18 : CLKBUF_X1 port map( A => n14, Z => n8);
   U19 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => n9);
   U20 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n69);
   U21 : NAND2_X2 port map( A1 => n11, A2 => n78, ZN => n99);
   U22 : BUF_X2 port map( A => n96, Z => n14);
   U23 : BUF_X1 port map( A => n94, Z => n12);
   U24 : BUF_X1 port map( A => n96, Z => n16);
   U25 : BUF_X1 port map( A => n98, Z => n17);
   U26 : BUF_X1 port map( A => n98, Z => n18);
   U27 : BUF_X1 port map( A => n98, Z => n19);
   U28 : INV_X1 port map( A => b(2), ZN => n61);
   U29 : INV_X1 port map( A => b(0), ZN => n24);
   U30 : INV_X1 port map( A => b(1), ZN => n78);
   U31 : NAND2_X1 port map( A1 => n2, A2 => n98, ZN => n23);
   U32 : XOR2_X1 port map( A => b(1), B => n10, Z => n21);
   U33 : NAND2_X1 port map( A1 => n21, A2 => n61, ZN => n94);
   U34 : MUX2_X1 port map( A => n23, B => n13, S => A(0), Z => n22);
   U35 : OAI211_X1 port map( C1 => n61, C2 => n85, A => n93, B => n22, ZN => 
                           p(0));
   U36 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n98);
   U37 : MUX2_X1 port map( A => n93, B => n19, S => A(0), Z => n26);
   U38 : NAND2_X1 port map( A1 => b(2), A2 => n69, ZN => n101);
   U39 : MUX2_X1 port map( A => n84, B => n13, S => A(1), Z => n25);
   U40 : NAND3_X1 port map( A1 => n26, A2 => n8, A3 => n25, ZN => p(1));
   U41 : MUX2_X1 port map( A => n93, B => n19, S => A(1), Z => n28);
   U42 : MUX2_X1 port map( A => n84, B => n13, S => A(2), Z => n27);
   U43 : NAND3_X1 port map( A1 => n28, A2 => n16, A3 => n27, ZN => p(2));
   U44 : MUX2_X1 port map( A => n99, B => n19, S => A(2), Z => n30);
   U45 : MUX2_X1 port map( A => n20, B => n12, S => A(3), Z => n29);
   U46 : NAND3_X1 port map( A1 => n30, A2 => n16, A3 => n29, ZN => p(3));
   U47 : MUX2_X1 port map( A => n93, B => n19, S => A(3), Z => n32);
   U48 : MUX2_X1 port map( A => n20, B => n12, S => A(4), Z => n31);
   U49 : NAND3_X1 port map( A1 => n32, A2 => n16, A3 => n31, ZN => p(4));
   U50 : MUX2_X1 port map( A => n93, B => n19, S => A(4), Z => n34);
   U51 : MUX2_X1 port map( A => n84, B => n12, S => A(5), Z => n33);
   U52 : NAND3_X1 port map( A1 => n34, A2 => n16, A3 => n33, ZN => p(5));
   U53 : MUX2_X1 port map( A => n99, B => n18, S => A(5), Z => n36);
   U54 : MUX2_X1 port map( A => n20, B => n12, S => A(6), Z => n35);
   U55 : NAND3_X1 port map( A1 => n36, A2 => n16, A3 => n35, ZN => p(6));
   U56 : MUX2_X1 port map( A => n99, B => n18, S => A(6), Z => n38);
   U57 : MUX2_X1 port map( A => n20, B => n12, S => A(7), Z => n37);
   U58 : NAND3_X1 port map( A1 => n38, A2 => n16, A3 => n37, ZN => p(7));
   U59 : MUX2_X1 port map( A => n93, B => n18, S => A(7), Z => n40);
   U60 : MUX2_X1 port map( A => n20, B => n12, S => A(8), Z => n39);
   U61 : NAND3_X1 port map( A1 => n40, A2 => n15, A3 => n39, ZN => p(8));
   U62 : MUX2_X1 port map( A => n99, B => n18, S => A(8), Z => n42);
   U63 : MUX2_X1 port map( A => n20, B => n12, S => A(9), Z => n41);
   U64 : NAND3_X1 port map( A1 => n42, A2 => n15, A3 => n41, ZN => p(9));
   U65 : MUX2_X1 port map( A => n93, B => n18, S => A(9), Z => n44);
   U66 : MUX2_X1 port map( A => n20, B => n12, S => A(10), Z => n43);
   U67 : NAND3_X1 port map( A1 => n44, A2 => n15, A3 => n43, ZN => p(10));
   U68 : MUX2_X1 port map( A => n99, B => n18, S => A(10), Z => n46);
   U69 : MUX2_X1 port map( A => n20, B => n12, S => A(11), Z => n45);
   U70 : NAND3_X1 port map( A1 => n46, A2 => n15, A3 => n45, ZN => p(11));
   U71 : MUX2_X1 port map( A => n99, B => n18, S => A(11), Z => n48);
   U72 : MUX2_X1 port map( A => n20, B => n12, S => A(12), Z => n47);
   U73 : NAND3_X1 port map( A1 => n48, A2 => n15, A3 => n47, ZN => p(12));
   U74 : MUX2_X1 port map( A => n99, B => n18, S => A(12), Z => n50);
   U75 : MUX2_X1 port map( A => n20, B => n12, S => A(13), Z => n49);
   U76 : NAND3_X1 port map( A1 => n50, A2 => n15, A3 => n49, ZN => p(13));
   U77 : MUX2_X1 port map( A => n99, B => n18, S => A(13), Z => n52);
   U78 : MUX2_X1 port map( A => n20, B => n1, S => A(14), Z => n51);
   U79 : NAND3_X1 port map( A1 => n52, A2 => n15, A3 => n51, ZN => p(14));
   U80 : MUX2_X1 port map( A => n99, B => n18, S => A(14), Z => n54);
   U81 : MUX2_X1 port map( A => n20, B => n13, S => A(15), Z => n53);
   U82 : NAND3_X1 port map( A1 => n54, A2 => n15, A3 => n53, ZN => p(15));
   U83 : MUX2_X1 port map( A => n99, B => n18, S => A(15), Z => n56);
   U84 : MUX2_X1 port map( A => n20, B => n1, S => A(16), Z => n55);
   U85 : NAND3_X1 port map( A1 => n55, A2 => n15, A3 => n56, ZN => p(16));
   U86 : MUX2_X1 port map( A => n93, B => n17, S => A(16), Z => n58);
   U87 : MUX2_X1 port map( A => n20, B => n1, S => A(17), Z => n57);
   U88 : NAND3_X1 port map( A1 => n58, A2 => n15, A3 => n57, ZN => p(17));
   U89 : MUX2_X1 port map( A => n99, B => n17, S => A(17), Z => n60);
   U90 : MUX2_X1 port map( A => n20, B => n1, S => A(18), Z => n59);
   U91 : NAND3_X1 port map( A1 => n60, A2 => n15, A3 => n59, ZN => p(18));
   U92 : MUX2_X1 port map( A => n99, B => n17, S => A(18), Z => n64);
   U93 : XOR2_X1 port map( A => b(0), B => b(1), Z => n62);
   U94 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => n83);
   U95 : MUX2_X1 port map( A => n20, B => n9, S => A(19), Z => n63);
   U96 : NAND3_X1 port map( A1 => n64, A2 => n7, A3 => n63, ZN => p(19));
   U97 : MUX2_X1 port map( A => n93, B => n17, S => A(19), Z => n66);
   U98 : MUX2_X1 port map( A => n20, B => n1, S => A(20), Z => n65);
   U99 : NAND3_X1 port map( A1 => n66, A2 => n8, A3 => n65, ZN => p(20));
   U100 : MUX2_X1 port map( A => n93, B => n17, S => A(20), Z => n68);
   U101 : MUX2_X1 port map( A => n20, B => n1, S => A(21), Z => n67);
   U102 : NAND3_X1 port map( A1 => n68, A2 => n7, A3 => n67, ZN => p(21));
   U103 : MUX2_X1 port map( A => n99, B => n17, S => A(21), Z => n71);
   U104 : NAND2_X1 port map( A1 => b(2), A2 => n69, ZN => n84);
   U105 : MUX2_X1 port map( A => n84, B => n9, S => A(22), Z => n70);
   U106 : NAND3_X1 port map( A1 => n71, A2 => n70, A3 => n14, ZN => p(22));
   U107 : NAND2_X1 port map( A1 => n10, A2 => b(1), ZN => n85);
   U108 : MUX2_X1 port map( A => n86, B => n85, S => A(22), Z => n73);
   U109 : NAND3_X1 port map( A1 => n72, A2 => n73, A3 => n14, ZN => p(23));
   U110 : MUX2_X1 port map( A => n84, B => n9, S => A(24), Z => n75);
   U111 : MUX2_X1 port map( A => n86, B => n17, S => A(23), Z => n74);
   U112 : NAND3_X1 port map( A1 => n16, A2 => n75, A3 => n74, ZN => p(24));
   U113 : MUX2_X1 port map( A => n84, B => n9, S => A(25), Z => n77);
   U114 : MUX2_X1 port map( A => n93, B => n85, S => A(24), Z => n76);
   U115 : NAND3_X1 port map( A1 => n77, A2 => n14, A3 => n76, ZN => p(25));
   U116 : MUX2_X1 port map( A => n84, B => n9, S => A(26), Z => n80);
   U117 : NAND2_X1 port map( A1 => n11, A2 => n78, ZN => n86);
   U118 : MUX2_X1 port map( A => n86, B => n85, S => A(25), Z => n79);
   U119 : NAND3_X1 port map( A1 => n80, A2 => n14, A3 => n79, ZN => p(26));
   U120 : MUX2_X1 port map( A => n93, B => n85, S => A(26), Z => n82);
   U121 : MUX2_X1 port map( A => n84, B => n1, S => A(27), Z => n81);
   U122 : NAND3_X1 port map( A1 => n82, A2 => n15, A3 => n81, ZN => p(27));
   U123 : MUX2_X1 port map( A => n84, B => n83, S => A(28), Z => n88);
   U124 : MUX2_X1 port map( A => n86, B => n85, S => A(27), Z => n87);
   U125 : NAND3_X1 port map( A1 => n88, A2 => n87, A3 => n14, ZN => p(28));
   U126 : MUX2_X1 port map( A => n99, B => n17, S => A(28), Z => n90);
   U127 : MUX2_X1 port map( A => n20, B => n1, S => A(29), Z => n89);
   U128 : NAND3_X1 port map( A1 => n90, A2 => n8, A3 => n89, ZN => p(29));
   U129 : MUX2_X1 port map( A => n93, B => n17, S => A(29), Z => n92);
   U130 : MUX2_X1 port map( A => n20, B => n1, S => A(30), Z => n91);
   U131 : NAND3_X1 port map( A1 => n92, A2 => n8, A3 => n91, ZN => p(30));
   U132 : MUX2_X1 port map( A => n99, B => n17, S => A(30), Z => n97);
   U133 : MUX2_X1 port map( A => n20, B => n1, S => A(31), Z => n95);
   U134 : NAND3_X1 port map( A1 => n97, A2 => n15, A3 => n95, ZN => p(31));
   U135 : MUX2_X1 port map( A => n99, B => n17, S => A(31), Z => n100);
   U136 : NAND2_X1 port map( A1 => n20, A2 => n100, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_14 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_14;

architecture SYN_beh of ENC_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105 : std_logic;

begin
   
   U3 : NAND2_X2 port map( A1 => n27, A2 => n76, ZN => n99);
   U4 : BUF_X2 port map( A => n99, Z => n17);
   U5 : BUF_X1 port map( A => n99, Z => n19);
   U6 : BUF_X1 port map( A => n99, Z => n18);
   U7 : CLKBUF_X1 port map( A => b(1), Z => n7);
   U8 : CLKBUF_X1 port map( A => b(0), Z => n4);
   U9 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n31);
   U10 : NAND2_X1 port map( A1 => n4, A2 => n1, ZN => n2);
   U11 : NAND2_X1 port map( A1 => n29, A2 => n7, ZN => n3);
   U12 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => n71);
   U13 : INV_X1 port map( A => n7, ZN => n1);
   U14 : BUF_X1 port map( A => n101, Z => n21);
   U15 : CLKBUF_X1 port map( A => n101, Z => n12);
   U16 : BUF_X2 port map( A => n105, Z => n9);
   U17 : BUF_X1 port map( A => n105, Z => n26);
   U18 : BUF_X2 port map( A => n101, Z => n13);
   U19 : CLKBUF_X1 port map( A => n101, Z => n20);
   U20 : CLKBUF_X1 port map( A => n9, Z => n5);
   U21 : NAND2_X1 port map( A1 => n27, A2 => n76, ZN => n6);
   U22 : BUF_X1 port map( A => b(1), Z => n8);
   U23 : NAND2_X2 port map( A1 => n14, A2 => n66, ZN => n103);
   U24 : BUF_X2 port map( A => n105, Z => n10);
   U25 : CLKBUF_X1 port map( A => n87, Z => n11);
   U26 : CLKBUF_X1 port map( A => n101, Z => n22);
   U27 : INV_X1 port map( A => n15, ZN => n87);
   U28 : BUF_X1 port map( A => n84, Z => n24);
   U29 : BUF_X1 port map( A => n84, Z => n23);
   U30 : CLKBUF_X1 port map( A => n84, Z => n25);
   U31 : AND2_X1 port map( A1 => n29, A2 => b(2), ZN => n14);
   U32 : AND2_X1 port map( A1 => n31, A2 => b(2), ZN => n15);
   U33 : NAND2_X1 port map( A1 => n14, A2 => n66, ZN => n16);
   U34 : INV_X1 port map( A => b(2), ZN => n76);
   U35 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n84);
   U36 : INV_X1 port map( A => b(0), ZN => n29);
   U37 : INV_X1 port map( A => b(1), ZN => n66);
   U38 : NAND2_X1 port map( A1 => n14, A2 => n66, ZN => n94);
   U39 : NAND2_X1 port map( A1 => b(2), A2 => n84, ZN => n30);
   U40 : XOR2_X1 port map( A => b(0), B => n8, Z => n27);
   U41 : MUX2_X1 port map( A => n30, B => n17, S => A(0), Z => n28);
   U42 : OAI211_X1 port map( C1 => n76, C2 => n84, A => n94, B => n28, ZN => 
                           p(0));
   U43 : MUX2_X1 port map( A => n16, B => n25, S => A(0), Z => n33);
   U44 : NAND2_X1 port map( A1 => n15, A2 => n30, ZN => n101);
   U45 : NAND2_X1 port map( A1 => n31, A2 => b(2), ZN => n105);
   U46 : MUX2_X1 port map( A => n26, B => n99, S => A(1), Z => n32);
   U47 : NAND3_X1 port map( A1 => n33, A2 => n12, A3 => n32, ZN => p(1));
   U48 : MUX2_X1 port map( A => n94, B => n25, S => A(1), Z => n35);
   U49 : MUX2_X1 port map( A => n5, B => n18, S => A(2), Z => n34);
   U50 : NAND3_X1 port map( A1 => n35, A2 => n22, A3 => n34, ZN => p(2));
   U51 : MUX2_X1 port map( A => n16, B => n25, S => A(2), Z => n37);
   U52 : MUX2_X1 port map( A => n10, B => n17, S => A(3), Z => n36);
   U53 : NAND3_X1 port map( A1 => n37, A2 => n20, A3 => n36, ZN => p(3));
   U54 : MUX2_X1 port map( A => n94, B => n25, S => A(3), Z => n39);
   U55 : MUX2_X1 port map( A => n5, B => n18, S => A(4), Z => n38);
   U56 : NAND3_X1 port map( A1 => n39, A2 => n12, A3 => n38, ZN => p(4));
   U57 : MUX2_X1 port map( A => n16, B => n25, S => A(4), Z => n41);
   U58 : MUX2_X1 port map( A => n26, B => n19, S => A(5), Z => n40);
   U59 : NAND3_X1 port map( A1 => n41, A2 => n13, A3 => n40, ZN => p(5));
   U60 : MUX2_X1 port map( A => n94, B => n25, S => A(5), Z => n43);
   U61 : MUX2_X1 port map( A => n10, B => n17, S => A(6), Z => n42);
   U62 : NAND3_X1 port map( A1 => n43, A2 => n22, A3 => n42, ZN => p(6));
   U63 : MUX2_X1 port map( A => n16, B => n25, S => A(6), Z => n45);
   U64 : MUX2_X1 port map( A => n5, B => n17, S => A(7), Z => n44);
   U65 : NAND3_X1 port map( A1 => n45, A2 => n20, A3 => n44, ZN => p(7));
   U66 : MUX2_X1 port map( A => n94, B => n25, S => A(7), Z => n47);
   U67 : MUX2_X1 port map( A => n5, B => n17, S => A(8), Z => n46);
   U68 : NAND3_X1 port map( A1 => n46, A2 => n12, A3 => n47, ZN => p(8));
   U69 : MUX2_X1 port map( A => n16, B => n24, S => A(8), Z => n49);
   U70 : MUX2_X1 port map( A => n9, B => n19, S => A(9), Z => n48);
   U71 : NAND3_X1 port map( A1 => n49, A2 => n20, A3 => n48, ZN => p(9));
   U72 : MUX2_X1 port map( A => n94, B => n24, S => A(9), Z => n51);
   U73 : MUX2_X1 port map( A => n10, B => n17, S => A(10), Z => n50);
   U74 : NAND3_X1 port map( A1 => n51, A2 => n13, A3 => n50, ZN => p(10));
   U75 : MUX2_X1 port map( A => n16, B => n24, S => A(10), Z => n53);
   U76 : MUX2_X1 port map( A => n10, B => n18, S => A(11), Z => n52);
   U77 : NAND3_X1 port map( A1 => n53, A2 => n22, A3 => n52, ZN => p(11));
   U78 : MUX2_X1 port map( A => n94, B => n24, S => A(11), Z => n55);
   U79 : MUX2_X1 port map( A => n10, B => n99, S => A(12), Z => n54);
   U80 : NAND3_X1 port map( A1 => n55, A2 => n22, A3 => n54, ZN => p(12));
   U81 : MUX2_X1 port map( A => n16, B => n24, S => A(12), Z => n57);
   U82 : MUX2_X1 port map( A => n10, B => n99, S => A(13), Z => n56);
   U83 : NAND3_X1 port map( A1 => n57, A2 => n22, A3 => n56, ZN => p(13));
   U84 : MUX2_X1 port map( A => n94, B => n24, S => A(13), Z => n59);
   U85 : MUX2_X1 port map( A => n26, B => n99, S => A(14), Z => n58);
   U86 : NAND3_X1 port map( A1 => n59, A2 => n12, A3 => n58, ZN => p(14));
   U87 : MUX2_X1 port map( A => n16, B => n24, S => A(14), Z => n61);
   U88 : MUX2_X1 port map( A => n10, B => n99, S => A(15), Z => n60);
   U89 : NAND3_X1 port map( A1 => n61, A2 => n12, A3 => n60, ZN => p(15));
   U90 : MUX2_X1 port map( A => n94, B => n24, S => A(15), Z => n63);
   U91 : MUX2_X1 port map( A => n26, B => n6, S => A(16), Z => n62);
   U92 : NAND3_X1 port map( A1 => n63, A2 => n20, A3 => n62, ZN => p(16));
   U93 : MUX2_X1 port map( A => n11, B => n99, S => A(17), Z => n65);
   U94 : MUX2_X1 port map( A => n16, B => n24, S => A(16), Z => n64);
   U95 : NAND3_X1 port map( A1 => n65, A2 => n13, A3 => n64, ZN => p(17));
   U96 : MUX2_X1 port map( A => n103, B => n24, S => A(17), Z => n68);
   U97 : MUX2_X1 port map( A => n10, B => n99, S => A(18), Z => n67);
   U98 : NAND3_X1 port map( A1 => n68, A2 => n13, A3 => n67, ZN => p(18));
   U99 : MUX2_X1 port map( A => n26, B => n17, S => A(19), Z => n70);
   U100 : MUX2_X1 port map( A => n94, B => n24, S => A(18), Z => n69);
   U101 : NAND3_X1 port map( A1 => n70, A2 => n13, A3 => n69, ZN => p(19));
   U102 : MUX2_X1 port map( A => n16, B => n23, S => A(19), Z => n73);
   U103 : NAND2_X1 port map( A1 => n71, A2 => n76, ZN => n81);
   U104 : MUX2_X1 port map( A => n9, B => n81, S => A(20), Z => n72);
   U105 : NAND3_X1 port map( A1 => n72, A2 => n21, A3 => n73, ZN => p(20));
   U106 : MUX2_X1 port map( A => n103, B => n23, S => A(20), Z => n75);
   U107 : MUX2_X1 port map( A => n9, B => n6, S => A(21), Z => n74);
   U108 : NAND3_X1 port map( A1 => n75, A2 => n13, A3 => n74, ZN => p(21));
   U109 : MUX2_X1 port map( A => n87, B => n81, S => A(22), Z => n78);
   U110 : MUX2_X1 port map( A => n103, B => n23, S => A(21), Z => n77);
   U111 : NAND3_X1 port map( A1 => n78, A2 => n13, A3 => n77, ZN => p(22));
   U112 : MUX2_X1 port map( A => n87, B => n81, S => A(23), Z => n80);
   U113 : MUX2_X1 port map( A => n103, B => n23, S => A(22), Z => n79);
   U114 : NAND3_X1 port map( A1 => n80, A2 => n79, A3 => n21, ZN => p(23));
   U115 : MUX2_X1 port map( A => n87, B => n81, S => A(24), Z => n83);
   U116 : MUX2_X1 port map( A => n103, B => n84, S => A(23), Z => n82);
   U117 : NAND3_X1 port map( A1 => n83, A2 => n21, A3 => n82, ZN => p(24));
   U118 : MUX2_X1 port map( A => n103, B => n84, S => A(24), Z => n86);
   U119 : MUX2_X1 port map( A => n87, B => n99, S => A(25), Z => n85);
   U120 : NAND3_X1 port map( A1 => n86, A2 => n13, A3 => n85, ZN => p(25));
   U121 : MUX2_X1 port map( A => n103, B => n23, S => A(25), Z => n89);
   U122 : MUX2_X1 port map( A => n11, B => n17, S => A(26), Z => n88);
   U123 : NAND3_X1 port map( A1 => n89, A2 => n88, A3 => n13, ZN => p(26));
   U124 : MUX2_X1 port map( A => n103, B => n23, S => A(26), Z => n91);
   U125 : MUX2_X1 port map( A => n10, B => n19, S => A(27), Z => n90);
   U126 : NAND3_X1 port map( A1 => n90, A2 => n21, A3 => n91, ZN => p(27));
   U127 : MUX2_X1 port map( A => n94, B => n23, S => A(27), Z => n93);
   U128 : MUX2_X1 port map( A => n26, B => n17, S => A(28), Z => n92);
   U129 : NAND3_X1 port map( A1 => n93, A2 => n92, A3 => n20, ZN => p(28));
   U130 : MUX2_X1 port map( A => n16, B => n23, S => A(28), Z => n96);
   U131 : MUX2_X1 port map( A => n10, B => n17, S => A(29), Z => n95);
   U132 : NAND3_X1 port map( A1 => n96, A2 => n13, A3 => n95, ZN => p(29));
   U133 : MUX2_X1 port map( A => n103, B => n23, S => A(29), Z => n98);
   U134 : MUX2_X1 port map( A => n9, B => n17, S => A(30), Z => n97);
   U135 : NAND3_X1 port map( A1 => n98, A2 => n13, A3 => n97, ZN => p(30));
   U136 : MUX2_X1 port map( A => n103, B => n23, S => A(30), Z => n102);
   U137 : MUX2_X1 port map( A => n9, B => n18, S => A(31), Z => n100);
   U138 : NAND3_X1 port map( A1 => n102, A2 => n12, A3 => n100, ZN => p(31));
   U139 : MUX2_X1 port map( A => n103, B => n23, S => A(31), Z => n104);
   U140 : NAND2_X1 port map( A1 => n9, A2 => n104, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_13 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_13;

architecture SYN_beh of ENC_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net29998, net30001, net30010, net30021, net30022, net30033, net30075,
      net30077, net30078, net30721, net31223, net31221, net31233, net31231, 
      net31227, net31424, net33597, net34021, net34028, net34047, net34495, 
      net34811, net36460, net37647, net37654, net37672, net37847, net42472, 
      net42478, net30030, net33339, net31219, n1, n2, n3, n4, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74 : std_logic;

begin
   
   U3 : BUF_X2 port map( A => n72, Z => n3);
   U4 : INV_X1 port map( A => net33339, ZN => net31219);
   U5 : AND3_X2 port map( A1 => n1, A2 => net30078, A3 => b(2), ZN => net33339)
                           ;
   U6 : MUX2_X1 port map( A => net31219, B => net34021, S => A(20), Z => 
                           net30030);
   U7 : MUX2_X1 port map( A => net31219, B => net34021, S => A(22), Z => 
                           net30022);
   U8 : INV_X1 port map( A => b(0), ZN => n1);
   U9 : INV_X1 port map( A => b(1), ZN => net30078);
   U10 : INV_X1 port map( A => net33339, ZN => net31221);
   U11 : INV_X1 port map( A => net33339, ZN => net34047);
   U12 : BUF_X1 port map( A => net33339, Z => net37647);
   U13 : NAND3_X1 port map( A1 => net30030, A2 => n2, A3 => net42472, ZN => 
                           p(21));
   U14 : CLKBUF_X1 port map( A => net30001, Z => net34021);
   U15 : MUX2_X1 port map( A => net30010, B => net29998, S => net30721, Z => n2
                           );
   U16 : NAND2_X1 port map( A1 => net33597, A2 => net30033, ZN => net30010);
   U17 : NAND2_X1 port map( A1 => net30075, A2 => net37847, ZN => net29998);
   U18 : INV_X1 port map( A => A(21), ZN => net30721);
   U19 : NAND2_X1 port map( A1 => net34028, A2 => net30077, ZN => net42472);
   U20 : CLKBUF_X1 port map( A => n72, Z => n4);
   U21 : BUF_X1 port map( A => net42472, Z => net31424);
   U22 : BUF_X1 port map( A => net42472, Z => net34495);
   U23 : CLKBUF_X1 port map( A => b(2), Z => net42478);
   U24 : INV_X1 port map( A => net31233, ZN => net31227);
   U25 : INV_X2 port map( A => net34028, ZN => net30021);
   U26 : INV_X2 port map( A => net31233, ZN => net31231);
   U27 : CLKBUF_X1 port map( A => b(2), Z => net37847);
   U28 : BUF_X1 port map( A => net29998, Z => net37672);
   U29 : INV_X1 port map( A => net29998, ZN => net37654);
   U30 : AND2_X1 port map( A1 => net30075, A2 => b(2), ZN => net34028);
   U31 : AND2_X1 port map( A1 => net37654, A2 => net30077, ZN => n5);
   U32 : INV_X1 port map( A => net37654, ZN => net36460);
   U33 : CLKBUF_X1 port map( A => b(1), Z => net34811);
   U34 : AND2_X1 port map( A1 => net37647, A2 => net30721, ZN => n6);
   U35 : AND2_X1 port map( A1 => A(21), A2 => net31233, ZN => n7);
   U36 : NOR3_X1 port map( A1 => n6, A2 => n7, A3 => n5, ZN => n54);
   U37 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => net30075);
   U38 : XNOR2_X1 port map( A => b(0), B => net30078, ZN => n8);
   U39 : XNOR2_X1 port map( A => b(0), B => net30078, ZN => net33597);
   U40 : INV_X1 port map( A => net30001, ZN => net31233);
   U41 : NAND2_X1 port map( A1 => n8, A2 => net30033, ZN => n9);
   U42 : INV_X1 port map( A => n5, ZN => n10);
   U43 : INV_X1 port map( A => net37647, ZN => net31223);
   U44 : INV_X1 port map( A => b(2), ZN => net30033);
   U45 : NAND2_X1 port map( A1 => net42478, A2 => net30001, ZN => net30077);
   U46 : NAND2_X1 port map( A1 => n8, A2 => net30033, ZN => n70);
   U47 : MUX2_X1 port map( A => net30077, B => n70, S => A(0), Z => n11);
   U48 : OAI211_X1 port map( C1 => net30033, C2 => net31231, A => net31223, B 
                           => n11, ZN => p(0));
   U49 : NAND2_X1 port map( A1 => b(0), A2 => net34811, ZN => net30001);
   U50 : MUX2_X1 port map( A => net31221, B => net31231, S => A(0), Z => n13);
   U51 : NAND2_X1 port map( A1 => net34028, A2 => net30077, ZN => n72);
   U52 : MUX2_X1 port map( A => net36460, B => n70, S => A(1), Z => n12);
   U53 : NAND3_X1 port map( A1 => n13, A2 => net31424, A3 => n12, ZN => p(1));
   U54 : MUX2_X1 port map( A => net31221, B => net31231, S => A(1), Z => n15);
   U55 : MUX2_X1 port map( A => net36460, B => n70, S => A(2), Z => n14);
   U56 : NAND3_X1 port map( A1 => n15, A2 => n10, A3 => n14, ZN => p(2));
   U57 : MUX2_X1 port map( A => net34047, B => net31231, S => A(2), Z => n17);
   U58 : MUX2_X1 port map( A => net36460, B => n70, S => A(3), Z => n16);
   U59 : NAND3_X1 port map( A1 => n17, A2 => n10, A3 => n16, ZN => p(3));
   U60 : MUX2_X1 port map( A => net34047, B => net31231, S => A(3), Z => n19);
   U61 : MUX2_X1 port map( A => net36460, B => n70, S => A(4), Z => n18);
   U62 : NAND3_X1 port map( A1 => n19, A2 => n10, A3 => n18, ZN => p(4));
   U63 : MUX2_X1 port map( A => net31221, B => net31231, S => A(4), Z => n21);
   U64 : MUX2_X1 port map( A => net36460, B => n9, S => A(5), Z => n20);
   U65 : NAND3_X1 port map( A1 => n21, A2 => n10, A3 => n20, ZN => p(5));
   U66 : MUX2_X1 port map( A => net31221, B => net31231, S => A(5), Z => n23);
   U67 : MUX2_X1 port map( A => net36460, B => n70, S => A(6), Z => n22);
   U68 : NAND3_X1 port map( A1 => n23, A2 => n10, A3 => n22, ZN => p(6));
   U69 : MUX2_X1 port map( A => net31221, B => net31231, S => A(6), Z => n25);
   U70 : MUX2_X1 port map( A => net36460, B => n9, S => A(7), Z => n24);
   U71 : NAND3_X1 port map( A1 => n25, A2 => n10, A3 => n24, ZN => p(7));
   U72 : MUX2_X1 port map( A => net34047, B => net31231, S => A(7), Z => n27);
   U73 : MUX2_X1 port map( A => net36460, B => n70, S => A(8), Z => n26);
   U74 : NAND3_X1 port map( A1 => n27, A2 => n3, A3 => n26, ZN => p(8));
   U75 : MUX2_X1 port map( A => net31223, B => net31231, S => A(8), Z => n29);
   U76 : MUX2_X1 port map( A => net36460, B => n70, S => A(9), Z => n28);
   U77 : NAND3_X1 port map( A1 => n29, A2 => net42472, A3 => n28, ZN => p(9));
   U78 : MUX2_X1 port map( A => net31221, B => net31231, S => A(9), Z => n31);
   U79 : MUX2_X1 port map( A => net30021, B => n9, S => A(10), Z => n30);
   U80 : NAND3_X1 port map( A1 => n31, A2 => net31424, A3 => n30, ZN => p(10));
   U81 : MUX2_X1 port map( A => net31221, B => net31231, S => A(10), Z => n33);
   U82 : MUX2_X1 port map( A => net30021, B => n70, S => A(11), Z => n32);
   U83 : NAND3_X1 port map( A1 => n33, A2 => net34495, A3 => n32, ZN => p(11));
   U84 : MUX2_X1 port map( A => net31223, B => net31231, S => A(11), Z => n35);
   U85 : MUX2_X1 port map( A => net30021, B => n9, S => A(12), Z => n34);
   U86 : NAND3_X1 port map( A1 => n35, A2 => net34495, A3 => n34, ZN => p(12));
   U87 : MUX2_X1 port map( A => net31223, B => net31231, S => A(12), Z => n37);
   U88 : MUX2_X1 port map( A => net30021, B => n70, S => A(13), Z => n36);
   U89 : NAND3_X1 port map( A1 => n37, A2 => net31424, A3 => n36, ZN => p(13));
   U90 : MUX2_X1 port map( A => net36460, B => n9, S => A(14), Z => n39);
   U91 : MUX2_X1 port map( A => net34047, B => net31231, S => A(13), Z => n38);
   U92 : NAND3_X1 port map( A1 => n39, A2 => n3, A3 => n38, ZN => p(14));
   U93 : MUX2_X1 port map( A => net37672, B => n50, S => A(15), Z => n41);
   U94 : MUX2_X1 port map( A => net34047, B => net31227, S => A(14), Z => n40);
   U95 : NAND3_X1 port map( A1 => n41, A2 => n3, A3 => n40, ZN => p(15));
   U96 : MUX2_X1 port map( A => net30021, B => n70, S => A(16), Z => n43);
   U97 : MUX2_X1 port map( A => net34047, B => net31231, S => A(15), Z => n42);
   U98 : NAND3_X1 port map( A1 => n43, A2 => n4, A3 => n42, ZN => p(16));
   U99 : MUX2_X1 port map( A => net30021, B => n9, S => A(17), Z => n45);
   U100 : MUX2_X1 port map( A => net31221, B => net31231, S => A(16), Z => n44)
                           ;
   U101 : NAND3_X1 port map( A1 => n45, A2 => net34495, A3 => n44, ZN => p(17))
                           ;
   U102 : MUX2_X1 port map( A => net31221, B => net31227, S => A(17), Z => n47)
                           ;
   U103 : NAND2_X1 port map( A1 => n8, A2 => net30033, ZN => n50);
   U104 : MUX2_X1 port map( A => net37672, B => n50, S => A(18), Z => n46);
   U105 : NAND3_X1 port map( A1 => n47, A2 => net34495, A3 => n46, ZN => p(18))
                           ;
   U106 : MUX2_X1 port map( A => net31221, B => net31227, S => A(18), Z => n49)
                           ;
   U107 : MUX2_X1 port map( A => net37672, B => n50, S => A(19), Z => n48);
   U108 : NAND3_X1 port map( A1 => n49, A2 => n4, A3 => n48, ZN => p(19));
   U109 : MUX2_X1 port map( A => net37672, B => n50, S => A(20), Z => n52);
   U110 : MUX2_X1 port map( A => net34047, B => net31227, S => A(19), Z => n51)
                           ;
   U111 : NAND3_X1 port map( A1 => n52, A2 => net31424, A3 => n51, ZN => p(20))
                           ;
   U112 : MUX2_X1 port map( A => net37672, B => n50, S => A(22), Z => n53);
   U113 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => p(22));
   U114 : MUX2_X1 port map( A => net29998, B => net30010, S => A(23), Z => n55)
                           ;
   U115 : NAND3_X1 port map( A1 => net30022, A2 => n55, A3 => net42472, ZN => 
                           p(23));
   U116 : MUX2_X1 port map( A => net34047, B => net31227, S => A(23), Z => n57)
                           ;
   U117 : MUX2_X1 port map( A => net37672, B => n9, S => A(24), Z => n56);
   U118 : NAND3_X1 port map( A1 => n57, A2 => n4, A3 => n56, ZN => p(24));
   U119 : MUX2_X1 port map( A => net31223, B => net31231, S => A(24), Z => n59)
                           ;
   U120 : MUX2_X1 port map( A => net30021, B => n9, S => A(25), Z => n58);
   U121 : NAND3_X1 port map( A1 => n59, A2 => net31424, A3 => n58, ZN => p(25))
                           ;
   U122 : MUX2_X1 port map( A => net34047, B => net31231, S => A(25), Z => n61)
                           ;
   U123 : MUX2_X1 port map( A => net36460, B => n9, S => A(26), Z => n60);
   U124 : NAND3_X1 port map( A1 => n61, A2 => n4, A3 => n60, ZN => p(26));
   U125 : MUX2_X1 port map( A => net36460, B => n9, S => A(27), Z => n63);
   U126 : MUX2_X1 port map( A => net31223, B => net31231, S => A(26), Z => n62)
                           ;
   U127 : NAND3_X1 port map( A1 => n63, A2 => n4, A3 => n62, ZN => p(27));
   U128 : MUX2_X1 port map( A => net31223, B => net31231, S => A(27), Z => n65)
                           ;
   U129 : MUX2_X1 port map( A => net30021, B => n9, S => A(28), Z => n64);
   U130 : NAND3_X1 port map( A1 => n65, A2 => n3, A3 => n64, ZN => p(28));
   U131 : MUX2_X1 port map( A => net30021, B => n50, S => A(29), Z => n67);
   U132 : MUX2_X1 port map( A => net34047, B => net31231, S => A(28), Z => n66)
                           ;
   U133 : NAND3_X1 port map( A1 => n67, A2 => n3, A3 => n66, ZN => p(29));
   U134 : MUX2_X1 port map( A => net31223, B => net31227, S => A(29), Z => n69)
                           ;
   U135 : MUX2_X1 port map( A => net30021, B => n50, S => A(30), Z => n68);
   U136 : NAND3_X1 port map( A1 => n69, A2 => net34495, A3 => n68, ZN => p(30))
                           ;
   U137 : MUX2_X1 port map( A => net31221, B => net31231, S => A(30), Z => n73)
                           ;
   U138 : MUX2_X1 port map( A => net30021, B => n9, S => A(31), Z => n71);
   U139 : NAND3_X1 port map( A1 => n73, A2 => n3, A3 => n71, ZN => p(31));
   U140 : MUX2_X1 port map( A => net34047, B => net31227, S => A(31), Z => n74)
                           ;
   U141 : NAND2_X1 port map( A1 => net30021, A2 => n74, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_12 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_12;

architecture SYN_beh of ENC_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net29919, net29922, net29924, net29927, net29930, net29949, net29954,
      net31195, net31193, net31201, net31199, net31197, net31207, net31203, 
      net31213, net31211, net31378, net31510, net31509, net31508, net31507, 
      net34050, net34049, net34150, net34191, net34266, net31205, net29996, 
      net29995, net29994, net29951, net29948, net29921, net37587, net34501, 
      net29964, net29952, net34310, net34125, net29926, n1, n2, n3, n4, n5, n6,
      n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63 : 
      std_logic;

begin
   
   U3 : CLKBUF_X1 port map( A => b(2), Z => n1);
   U4 : INV_X1 port map( A => b(1), ZN => n2);
   U5 : BUF_X1 port map( A => b(2), Z => net34310);
   U6 : BUF_X4 port map( A => net29921, Z => net31193);
   U7 : NAND2_X1 port map( A1 => net29964, A2 => net37587, ZN => net31213);
   U8 : NAND2_X1 port map( A1 => n3, A2 => net34310, ZN => net29926);
   U9 : MUX2_X1 port map( A => net29926, B => net34501, S => A(19), Z => 
                           net29952);
   U10 : NAND2_X1 port map( A1 => net34310, A2 => net34125, ZN => net29919);
   U11 : NAND2_X1 port map( A1 => net34310, A2 => net29994, ZN => net29924);
   U12 : NAND2_X1 port map( A1 => n3, A2 => net34310, ZN => net34191);
   U13 : NAND2_X1 port map( A1 => net31508, A2 => n2, ZN => n3);
   U14 : NAND2_X1 port map( A1 => n4, A2 => n2, ZN => net34125);
   U15 : NAND3_X1 port map( A1 => net31508, A2 => b(2), A3 => net31507, ZN => 
                           net29921);
   U16 : INV_X1 port map( A => b(0), ZN => n4);
   U17 : NAND2_X1 port map( A1 => net29995, A2 => n1, ZN => net29994);
   U18 : INV_X1 port map( A => b(2), ZN => net29964);
   U19 : NAND3_X1 port map( A1 => net29952, A2 => net29951, A3 => net31205, ZN 
                           => p(19));
   U20 : NAND2_X1 port map( A1 => n5, A2 => net29964, ZN => net34501);
   U21 : MUX2_X1 port map( A => net29919, B => net34501, S => A(21), Z => 
                           net29948);
   U22 : NAND2_X1 port map( A1 => net37587, A2 => net29964, ZN => net29930);
   U23 : OAI211_X1 port map( C1 => net29964, C2 => net31199, A => net31193, B 
                           => net29996, ZN => p(0));
   U24 : NAND2_X1 port map( A1 => net37587, A2 => net29964, ZN => net29927);
   U25 : NAND2_X1 port map( A1 => net31509, A2 => net31510, ZN => n5);
   U26 : MUX2_X1 port map( A => net31195, B => net31199, S => A(19), Z => 
                           net29949);
   U27 : NAND2_X1 port map( A1 => net31509, A2 => net31510, ZN => net37587);
   U28 : BUF_X1 port map( A => net29924, Z => net31205);
   U29 : NAND3_X1 port map( A1 => net29948, A2 => n6, A3 => net31205, ZN => 
                           p(21));
   U30 : MUX2_X1 port map( A => net29921, B => net29995, S => A(18), Z => 
                           net29951);
   U31 : CLKBUF_X1 port map( A => net29921, Z => net31195);
   U32 : MUX2_X1 port map( A => net29921, B => net31199, S => A(20), Z => n6);
   U33 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => net29995);
   U34 : MUX2_X1 port map( A => net34191, B => net29927, S => A(18), Z => 
                           net29954);
   U35 : MUX2_X1 port map( A => net29994, B => net31211, S => A(0), Z => 
                           net29996);
   U36 : CLKBUF_X1 port map( A => net29919, Z => net34150);
   U37 : BUF_X2 port map( A => net29922, Z => net31199);
   U38 : CLKBUF_X1 port map( A => net29927, Z => net31211);
   U39 : BUF_X1 port map( A => net29924, Z => net34266);
   U40 : BUF_X1 port map( A => net29924, Z => net34049);
   U41 : BUF_X1 port map( A => net29924, Z => net34050);
   U42 : BUF_X2 port map( A => net29919, Z => net31378);
   U43 : CLKBUF_X1 port map( A => net29922, Z => net31197);
   U44 : BUF_X1 port map( A => net29924, Z => net31203);
   U45 : CLKBUF_X1 port map( A => net29924, Z => net31207);
   U46 : CLKBUF_X1 port map( A => net29922, Z => net31201);
   U47 : NAND2_X1 port map( A1 => b(1), A2 => n4, ZN => net31509);
   U48 : NAND2_X1 port map( A1 => net31507, A2 => b(0), ZN => net31510);
   U49 : INV_X1 port map( A => b(1), ZN => net31507);
   U50 : INV_X1 port map( A => b(0), ZN => net31508);
   U51 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => net29922);
   U52 : MUX2_X1 port map( A => net31193, B => net31201, S => A(0), Z => n8);
   U53 : MUX2_X1 port map( A => net31378, B => net31211, S => A(1), Z => n7);
   U54 : NAND3_X1 port map( A1 => n8, A2 => net31203, A3 => n7, ZN => p(1));
   U55 : MUX2_X1 port map( A => net31193, B => net31201, S => A(1), Z => n10);
   U56 : MUX2_X1 port map( A => net31378, B => net31211, S => A(2), Z => n9);
   U57 : NAND3_X1 port map( A1 => n10, A2 => net34049, A3 => n9, ZN => p(2));
   U58 : MUX2_X1 port map( A => net31193, B => net31201, S => A(2), Z => n12);
   U59 : MUX2_X1 port map( A => net31378, B => net31211, S => A(3), Z => n11);
   U60 : NAND3_X1 port map( A1 => n12, A2 => net34050, A3 => n11, ZN => p(3));
   U61 : MUX2_X1 port map( A => net31193, B => net31201, S => A(3), Z => n14);
   U62 : MUX2_X1 port map( A => net31378, B => net31211, S => A(4), Z => n13);
   U63 : NAND3_X1 port map( A1 => n14, A2 => net31207, A3 => n13, ZN => p(4));
   U64 : MUX2_X1 port map( A => net31193, B => net31201, S => A(4), Z => n16);
   U65 : MUX2_X1 port map( A => net31378, B => net31211, S => A(5), Z => n15);
   U66 : NAND3_X1 port map( A1 => n16, A2 => net31203, A3 => n15, ZN => p(5));
   U67 : MUX2_X1 port map( A => net31193, B => net31201, S => A(5), Z => n18);
   U68 : MUX2_X1 port map( A => net31378, B => net31213, S => A(6), Z => n17);
   U69 : NAND3_X1 port map( A1 => n18, A2 => net31203, A3 => n17, ZN => p(6));
   U70 : MUX2_X1 port map( A => net31193, B => net31201, S => A(6), Z => n20);
   U71 : MUX2_X1 port map( A => net31378, B => net31213, S => A(7), Z => n19);
   U72 : NAND3_X1 port map( A1 => n20, A2 => net34266, A3 => n19, ZN => p(7));
   U73 : MUX2_X1 port map( A => net31193, B => net31201, S => A(7), Z => n22);
   U74 : MUX2_X1 port map( A => net31378, B => net29930, S => A(8), Z => n21);
   U75 : NAND3_X1 port map( A1 => n22, A2 => net31207, A3 => n21, ZN => p(8));
   U76 : MUX2_X1 port map( A => net31193, B => net31201, S => A(8), Z => n24);
   U77 : MUX2_X1 port map( A => net31378, B => net31213, S => A(9), Z => n23);
   U78 : NAND3_X1 port map( A1 => n24, A2 => net34049, A3 => n23, ZN => p(9));
   U79 : MUX2_X1 port map( A => net31193, B => net31201, S => A(9), Z => n26);
   U80 : MUX2_X1 port map( A => net34191, B => net29927, S => A(10), Z => n25);
   U81 : NAND3_X1 port map( A1 => n26, A2 => net31203, A3 => n25, ZN => p(10));
   U82 : MUX2_X1 port map( A => net31193, B => net31199, S => A(10), Z => n28);
   U83 : MUX2_X1 port map( A => net31378, B => net29930, S => A(11), Z => n27);
   U84 : NAND3_X1 port map( A1 => n28, A2 => net34266, A3 => n27, ZN => p(11));
   U85 : MUX2_X1 port map( A => net31193, B => net31199, S => A(11), Z => n30);
   U86 : MUX2_X1 port map( A => net34191, B => net29927, S => A(12), Z => n29);
   U87 : NAND3_X1 port map( A1 => n30, A2 => net34049, A3 => n29, ZN => p(12));
   U88 : MUX2_X1 port map( A => net31195, B => net31199, S => A(12), Z => n32);
   U89 : MUX2_X1 port map( A => net34150, B => net29930, S => A(13), Z => n31);
   U90 : NAND3_X1 port map( A1 => n32, A2 => net34049, A3 => n31, ZN => p(13));
   U91 : MUX2_X1 port map( A => net34191, B => net31213, S => A(14), Z => n34);
   U92 : MUX2_X1 port map( A => net31193, B => net31199, S => A(13), Z => n33);
   U93 : NAND3_X1 port map( A1 => n34, A2 => net34050, A3 => n33, ZN => p(14));
   U94 : MUX2_X1 port map( A => net31193, B => net31199, S => A(14), Z => n36);
   U95 : MUX2_X1 port map( A => net31378, B => net31213, S => A(15), Z => n35);
   U96 : NAND3_X1 port map( A1 => n36, A2 => net34049, A3 => n35, ZN => p(15));
   U97 : MUX2_X1 port map( A => net31193, B => net31199, S => A(15), Z => n38);
   U98 : MUX2_X1 port map( A => net34191, B => net29927, S => A(16), Z => n37);
   U99 : NAND3_X1 port map( A1 => n38, A2 => net31207, A3 => n37, ZN => p(16));
   U100 : MUX2_X1 port map( A => net31193, B => net31199, S => A(16), Z => n40)
                           ;
   U101 : MUX2_X1 port map( A => net31378, B => net29930, S => A(17), Z => n39)
                           ;
   U102 : NAND3_X1 port map( A1 => n40, A2 => net34266, A3 => n39, ZN => p(17))
                           ;
   U103 : MUX2_X1 port map( A => net31195, B => net31199, S => A(17), Z => n41)
                           ;
   U104 : NAND3_X1 port map( A1 => n41, A2 => net29954, A3 => net34050, ZN => 
                           p(18));
   U105 : MUX2_X1 port map( A => net34150, B => net29930, S => A(20), Z => n42)
                           ;
   U106 : NAND3_X1 port map( A1 => net29949, A2 => n42, A3 => net34266, ZN => 
                           p(20));
   U107 : MUX2_X1 port map( A => net31193, B => net31197, S => A(21), Z => n44)
                           ;
   U108 : MUX2_X1 port map( A => net34191, B => net29927, S => A(22), Z => n43)
                           ;
   U109 : NAND3_X1 port map( A1 => n44, A2 => net34266, A3 => n43, ZN => p(22))
                           ;
   U110 : MUX2_X1 port map( A => net31195, B => net31197, S => A(22), Z => n46)
                           ;
   U111 : MUX2_X1 port map( A => net34150, B => net29930, S => A(23), Z => n45)
                           ;
   U112 : NAND3_X1 port map( A1 => n46, A2 => net31203, A3 => n45, ZN => p(23))
                           ;
   U113 : MUX2_X1 port map( A => net31193, B => net31197, S => A(23), Z => n48)
                           ;
   U114 : MUX2_X1 port map( A => net34191, B => net31211, S => A(24), Z => n47)
                           ;
   U115 : NAND3_X1 port map( A1 => n48, A2 => net31207, A3 => n47, ZN => p(24))
                           ;
   U116 : MUX2_X1 port map( A => net31193, B => net31197, S => A(24), Z => n50)
                           ;
   U117 : MUX2_X1 port map( A => net31378, B => net31211, S => A(25), Z => n49)
                           ;
   U118 : NAND3_X1 port map( A1 => n50, A2 => net34266, A3 => n49, ZN => p(25))
                           ;
   U119 : MUX2_X1 port map( A => net31193, B => net31197, S => A(25), Z => n52)
                           ;
   U120 : MUX2_X1 port map( A => net31378, B => net29927, S => A(26), Z => n51)
                           ;
   U121 : NAND3_X1 port map( A1 => n52, A2 => net31203, A3 => n51, ZN => p(26))
                           ;
   U122 : MUX2_X1 port map( A => net31193, B => net31197, S => A(26), Z => n54)
                           ;
   U123 : MUX2_X1 port map( A => net31378, B => net29927, S => A(27), Z => n53)
                           ;
   U124 : NAND3_X1 port map( A1 => n54, A2 => net34266, A3 => n53, ZN => p(27))
                           ;
   U125 : MUX2_X1 port map( A => net31195, B => net31197, S => A(27), Z => n56)
                           ;
   U126 : MUX2_X1 port map( A => net34191, B => net31211, S => A(28), Z => n55)
                           ;
   U127 : NAND3_X1 port map( A1 => n56, A2 => net34050, A3 => n55, ZN => p(28))
                           ;
   U128 : MUX2_X1 port map( A => net31193, B => net31197, S => A(28), Z => n58)
                           ;
   U129 : MUX2_X1 port map( A => net34191, B => net31211, S => A(29), Z => n57)
                           ;
   U130 : NAND3_X1 port map( A1 => n58, A2 => net34049, A3 => n57, ZN => p(29))
                           ;
   U131 : MUX2_X1 port map( A => net31193, B => net31197, S => A(29), Z => n60)
                           ;
   U132 : MUX2_X1 port map( A => net31378, B => net31211, S => A(30), Z => n59)
                           ;
   U133 : NAND3_X1 port map( A1 => n60, A2 => net34050, A3 => n59, ZN => p(30))
                           ;
   U134 : MUX2_X1 port map( A => net31193, B => net31197, S => A(30), Z => n62)
                           ;
   U135 : MUX2_X1 port map( A => net34191, B => net31211, S => A(31), Z => n61)
                           ;
   U136 : NAND3_X1 port map( A1 => n62, A2 => net34050, A3 => n61, ZN => p(31))
                           ;
   U137 : MUX2_X1 port map( A => net31195, B => net31197, S => A(31), Z => n63)
                           ;
   U138 : NAND2_X1 port map( A1 => net31378, A2 => n63, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_11 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_11;

architecture SYN_beh of ENC_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n33, A2 => n15, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n32, A2 => n34, ZN => n2);
   U5 : AND3_X1 port map( A1 => n1, A2 => n2, A3 => n25, ZN => n86);
   U6 : NAND3_X1 port map( A1 => n14, A2 => n58, A3 => n59, ZN => p(11));
   U7 : CLKBUF_X1 port map( A => b(0), Z => n3);
   U8 : CLKBUF_X1 port map( A => n72, Z => n4);
   U9 : CLKBUF_X1 port map( A => n73, Z => n28);
   U10 : BUF_X2 port map( A => n73, Z => n27);
   U11 : NAND2_X1 port map( A1 => n18, A2 => n8, ZN => n102);
   U12 : NAND2_X1 port map( A1 => n19, A2 => n79, ZN => n5);
   U13 : AND2_X1 port map( A1 => n7, A2 => n79, ZN => n6);
   U14 : INV_X1 port map( A => n17, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n7);
   U16 : INV_X2 port map( A => n15, ZN => n20);
   U17 : NAND2_X1 port map( A1 => b(0), A2 => n8, ZN => n9);
   U18 : NAND2_X1 port map( A1 => n35, A2 => b(1), ZN => n10);
   U19 : NAND2_X1 port map( A1 => n10, A2 => n9, ZN => n19);
   U20 : INV_X1 port map( A => b(1), ZN => n8);
   U21 : CLKBUF_X1 port map( A => n16, Z => n11);
   U22 : CLKBUF_X1 port map( A => n31, Z => n12);
   U23 : INV_X1 port map( A => n17, ZN => n13);
   U24 : INV_X1 port map( A => n17, ZN => n14);
   U25 : INV_X1 port map( A => n17, ZN => n23);
   U26 : INV_X1 port map( A => n97, ZN => n15);
   U27 : INV_X1 port map( A => n32, ZN => n16);
   U28 : INV_X1 port map( A => n32, ZN => n31);
   U29 : CLKBUF_X1 port map( A => n73, Z => n26);
   U30 : BUF_X2 port map( A => n110, Z => n29);
   U31 : BUF_X2 port map( A => n102, Z => n30);
   U32 : AND2_X2 port map( A1 => n37, A2 => n72, ZN => n17);
   U33 : AND2_X1 port map( A1 => b(2), A2 => n35, ZN => n18);
   U34 : INV_X1 port map( A => n6, ZN => n21);
   U35 : INV_X1 port map( A => n6, ZN => n22);
   U36 : INV_X1 port map( A => n17, ZN => n25);
   U37 : INV_X1 port map( A => n112, ZN => n32);
   U38 : INV_X1 port map( A => n34, ZN => n33);
   U39 : INV_X1 port map( A => A(21), ZN => n34);
   U40 : INV_X1 port map( A => b(2), ZN => n79);
   U41 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n73);
   U42 : INV_X1 port map( A => b(0), ZN => n35);
   U43 : NAND2_X1 port map( A1 => n18, A2 => n8, ZN => n110);
   U44 : NAND2_X1 port map( A1 => b(2), A2 => n73, ZN => n72);
   U45 : NAND2_X1 port map( A1 => n19, A2 => n79, ZN => n107);
   U46 : MUX2_X1 port map( A => n4, B => n20, S => A(0), Z => n36);
   U47 : OAI211_X1 port map( C1 => n79, C2 => n28, A => n29, B => n36, ZN => 
                           p(0));
   U48 : MUX2_X1 port map( A => n29, B => n28, S => A(0), Z => n39);
   U49 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => b(2), ZN => n82);
   U50 : INV_X1 port map( A => n82, ZN => n37);
   U51 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => b(2), ZN => n112);
   U52 : MUX2_X1 port map( A => n31, B => n20, S => A(1), Z => n38);
   U53 : NAND3_X1 port map( A1 => n39, A2 => n24, A3 => n38, ZN => p(1));
   U54 : MUX2_X1 port map( A => n29, B => n28, S => A(1), Z => n41);
   U55 : MUX2_X1 port map( A => n16, B => n20, S => A(2), Z => n40);
   U56 : NAND3_X1 port map( A1 => n41, A2 => n13, A3 => n40, ZN => p(2));
   U57 : MUX2_X1 port map( A => n29, B => n28, S => A(2), Z => n43);
   U58 : MUX2_X1 port map( A => n11, B => n20, S => A(3), Z => n42);
   U59 : NAND3_X1 port map( A1 => n43, A2 => n14, A3 => n42, ZN => p(3));
   U60 : MUX2_X1 port map( A => n29, B => n28, S => A(3), Z => n45);
   U61 : MUX2_X1 port map( A => n11, B => n21, S => A(4), Z => n44);
   U62 : NAND3_X1 port map( A1 => n45, A2 => n24, A3 => n44, ZN => p(4));
   U63 : MUX2_X1 port map( A => n29, B => n28, S => A(4), Z => n47);
   U64 : MUX2_X1 port map( A => n16, B => n20, S => A(5), Z => n46);
   U65 : NAND3_X1 port map( A1 => n47, A2 => n24, A3 => n46, ZN => p(5));
   U66 : MUX2_X1 port map( A => n29, B => n28, S => A(5), Z => n49);
   U67 : MUX2_X1 port map( A => n16, B => n20, S => A(6), Z => n48);
   U68 : NAND3_X1 port map( A1 => n49, A2 => n23, A3 => n48, ZN => p(6));
   U69 : MUX2_X1 port map( A => n29, B => n28, S => A(6), Z => n51);
   U70 : MUX2_X1 port map( A => n12, B => n20, S => A(7), Z => n50);
   U71 : NAND3_X1 port map( A1 => n51, A2 => n23, A3 => n50, ZN => p(7));
   U72 : MUX2_X1 port map( A => n29, B => n28, S => A(7), Z => n53);
   U73 : MUX2_X1 port map( A => n31, B => n21, S => A(8), Z => n52);
   U74 : NAND3_X1 port map( A1 => n53, A2 => n14, A3 => n52, ZN => p(8));
   U75 : MUX2_X1 port map( A => n29, B => n28, S => A(8), Z => n55);
   U76 : MUX2_X1 port map( A => n11, B => n21, S => A(9), Z => n54);
   U77 : NAND3_X1 port map( A1 => n55, A2 => n14, A3 => n54, ZN => p(9));
   U78 : MUX2_X1 port map( A => n31, B => n20, S => A(10), Z => n57);
   U79 : MUX2_X1 port map( A => n29, B => n27, S => A(9), Z => n56);
   U80 : NAND3_X1 port map( A1 => n57, A2 => n13, A3 => n56, ZN => p(10));
   U81 : MUX2_X1 port map( A => n29, B => n27, S => A(10), Z => n59);
   U82 : MUX2_X1 port map( A => n31, B => n20, S => A(11), Z => n58);
   U83 : MUX2_X1 port map( A => n29, B => n27, S => A(11), Z => n61);
   U84 : MUX2_X1 port map( A => n31, B => n22, S => A(12), Z => n60);
   U85 : NAND3_X1 port map( A1 => n61, A2 => n24, A3 => n60, ZN => p(12));
   U86 : MUX2_X1 port map( A => n29, B => n27, S => A(12), Z => n63);
   U87 : MUX2_X1 port map( A => n16, B => n20, S => A(13), Z => n62);
   U88 : NAND3_X1 port map( A1 => n63, A2 => n23, A3 => n62, ZN => p(13));
   U89 : MUX2_X1 port map( A => n29, B => n27, S => A(13), Z => n65);
   U90 : MUX2_X1 port map( A => n11, B => n21, S => A(14), Z => n64);
   U91 : NAND3_X1 port map( A1 => n65, A2 => n23, A3 => n64, ZN => p(14));
   U92 : MUX2_X1 port map( A => n30, B => n27, S => A(14), Z => n67);
   U93 : MUX2_X1 port map( A => n11, B => n21, S => A(15), Z => n66);
   U94 : NAND3_X1 port map( A1 => n67, A2 => n23, A3 => n66, ZN => p(15));
   U95 : MUX2_X1 port map( A => n110, B => n27, S => A(15), Z => n69);
   U96 : NAND2_X1 port map( A1 => n7, A2 => n79, ZN => n97);
   U97 : MUX2_X1 port map( A => n31, B => n5, S => A(16), Z => n68);
   U98 : NAND3_X1 port map( A1 => n69, A2 => n23, A3 => n68, ZN => p(16));
   U99 : MUX2_X1 port map( A => n110, B => n27, S => A(16), Z => n71);
   U100 : MUX2_X1 port map( A => n31, B => n5, S => A(17), Z => n70);
   U101 : NAND3_X1 port map( A1 => n71, A2 => n13, A3 => n70, ZN => p(17));
   U102 : INV_X1 port map( A => n4, ZN => n76);
   U103 : MUX2_X1 port map( A => n102, B => n73, S => A(17), Z => n75);
   U104 : MUX2_X1 port map( A => n82, B => n107, S => A(18), Z => n74);
   U105 : OAI211_X1 port map( C1 => n76, C2 => n82, A => n75, B => n74, ZN => 
                           p(18));
   U106 : MUX2_X1 port map( A => n82, B => n97, S => A(19), Z => n78);
   U107 : MUX2_X1 port map( A => n102, B => n27, S => A(18), Z => n77);
   U108 : NAND3_X1 port map( A1 => n25, A2 => n78, A3 => n77, ZN => p(19));
   U109 : XOR2_X1 port map( A => b(1), B => n3, Z => n80);
   U110 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => n81);
   U111 : MUX2_X1 port map( A => n82, B => n81, S => A(20), Z => n84);
   U112 : MUX2_X1 port map( A => n110, B => n27, S => A(19), Z => n83);
   U113 : NAND3_X1 port map( A1 => n84, A2 => n23, A3 => n83, ZN => p(20));
   U114 : MUX2_X1 port map( A => n30, B => n27, S => A(20), Z => n85);
   U115 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => p(21));
   U116 : MUX2_X1 port map( A => n110, B => n26, S => n33, Z => n88);
   U117 : MUX2_X1 port map( A => n16, B => n5, S => A(22), Z => n87);
   U118 : NAND3_X1 port map( A1 => n88, A2 => n24, A3 => n87, ZN => p(22));
   U119 : MUX2_X1 port map( A => n16, B => n22, S => A(23), Z => n90);
   U120 : MUX2_X1 port map( A => n30, B => n26, S => A(22), Z => n89);
   U121 : NAND3_X1 port map( A1 => n90, A2 => n13, A3 => n89, ZN => p(23));
   U122 : MUX2_X1 port map( A => n30, B => n26, S => A(23), Z => n92);
   U123 : MUX2_X1 port map( A => n12, B => n21, S => A(24), Z => n91);
   U124 : NAND3_X1 port map( A1 => n92, A2 => n13, A3 => n91, ZN => p(24));
   U125 : MUX2_X1 port map( A => n30, B => n26, S => A(24), Z => n94);
   U126 : MUX2_X1 port map( A => n31, B => n21, S => A(25), Z => n93);
   U127 : NAND3_X1 port map( A1 => n94, A2 => n24, A3 => n93, ZN => p(25));
   U128 : MUX2_X1 port map( A => n16, B => n5, S => A(26), Z => n96);
   U129 : MUX2_X1 port map( A => n30, B => n26, S => A(25), Z => n95);
   U130 : NAND3_X1 port map( A1 => n96, A2 => n13, A3 => n95, ZN => p(26));
   U131 : MUX2_X1 port map( A => n110, B => n26, S => A(26), Z => n99);
   U132 : MUX2_X1 port map( A => n112, B => n5, S => A(27), Z => n98);
   U133 : NAND3_X1 port map( A1 => n99, A2 => n25, A3 => n98, ZN => p(27));
   U134 : MUX2_X1 port map( A => n30, B => n26, S => A(27), Z => n101);
   U135 : MUX2_X1 port map( A => n16, B => n21, S => A(28), Z => n100);
   U136 : NAND3_X1 port map( A1 => n101, A2 => n14, A3 => n100, ZN => p(28));
   U137 : MUX2_X1 port map( A => n110, B => n26, S => A(28), Z => n104);
   U138 : MUX2_X1 port map( A => n31, B => n21, S => A(29), Z => n103);
   U139 : NAND3_X1 port map( A1 => n104, A2 => n14, A3 => n103, ZN => p(29));
   U140 : MUX2_X1 port map( A => n30, B => n26, S => A(29), Z => n106);
   U141 : MUX2_X1 port map( A => n16, B => n20, S => A(30), Z => n105);
   U142 : NAND3_X1 port map( A1 => n106, A2 => n24, A3 => n105, ZN => p(30));
   U143 : MUX2_X1 port map( A => n30, B => n26, S => A(30), Z => n109);
   U144 : MUX2_X1 port map( A => n31, B => n21, S => A(31), Z => n108);
   U145 : NAND3_X1 port map( A1 => n109, A2 => n14, A3 => n108, ZN => p(31));
   U146 : MUX2_X1 port map( A => n30, B => n26, S => A(31), Z => n111);
   U147 : NAND2_X1 port map( A1 => n12, A2 => n111, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_10 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_10;

architecture SYN_beh of ENC_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96 : std_logic;

begin
   
   U3 : NAND2_X2 port map( A1 => n60, A2 => n5, ZN => n18);
   U4 : AND2_X2 port map( A1 => b(2), A2 => n22, ZN => n5);
   U5 : CLKBUF_X3 port map( A => n94, Z => n17);
   U6 : BUF_X2 port map( A => n76, Z => n9);
   U7 : BUF_X2 port map( A => n96, Z => n19);
   U8 : NAND2_X1 port map( A1 => b(0), A2 => n2, ZN => n3);
   U9 : NAND2_X1 port map( A1 => n1, A2 => b(1), ZN => n4);
   U10 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n6);
   U11 : INV_X1 port map( A => b(0), ZN => n1);
   U12 : INV_X1 port map( A => b(1), ZN => n2);
   U13 : BUF_X2 port map( A => n91, Z => n11);
   U14 : BUF_X2 port map( A => n96, Z => n21);
   U15 : BUF_X2 port map( A => n76, Z => n8);
   U16 : CLKBUF_X1 port map( A => n93, Z => n14);
   U17 : CLKBUF_X1 port map( A => n93, Z => n16);
   U18 : CLKBUF_X1 port map( A => n89, Z => n10);
   U19 : BUF_X2 port map( A => n91, Z => n12);
   U20 : BUF_X2 port map( A => n96, Z => n20);
   U21 : BUF_X1 port map( A => n93, Z => n15);
   U22 : BUF_X1 port map( A => n91, Z => n13);
   U23 : INV_X1 port map( A => n22, ZN => n7);
   U24 : NAND3_X1 port map( A1 => b(1), A2 => n7, A3 => b(2), ZN => n24);
   U25 : INV_X1 port map( A => b(0), ZN => n22);
   U26 : INV_X1 port map( A => b(1), ZN => n60);
   U27 : NAND2_X1 port map( A1 => n5, A2 => n60, ZN => n94);
   U28 : INV_X1 port map( A => b(2), ZN => n43);
   U29 : NAND2_X1 port map( A1 => n6, A2 => n43, ZN => n89);
   U30 : MUX2_X1 port map( A => n43, B => n10, S => A(0), Z => n23);
   U31 : NAND3_X1 port map( A1 => n24, A2 => n17, A3 => n23, ZN => p(0));
   U32 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n93);
   U33 : MUX2_X1 port map( A => n17, B => n16, S => A(0), Z => n26);
   U34 : NAND3_X1 port map( A1 => n7, A2 => b(2), A3 => b(1), ZN => n91);
   U35 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => b(2), ZN => n96);
   U36 : MUX2_X1 port map( A => n19, B => n10, S => A(1), Z => n25);
   U37 : NAND3_X1 port map( A1 => n26, A2 => n11, A3 => n25, ZN => p(1));
   U38 : MUX2_X1 port map( A => n17, B => n16, S => A(1), Z => n28);
   U39 : MUX2_X1 port map( A => n20, B => n9, S => A(2), Z => n27);
   U40 : NAND3_X1 port map( A1 => n28, A2 => n13, A3 => n27, ZN => p(2));
   U41 : MUX2_X1 port map( A => n17, B => n16, S => A(2), Z => n30);
   U42 : MUX2_X1 port map( A => n19, B => n9, S => A(3), Z => n29);
   U43 : NAND3_X1 port map( A1 => n30, A2 => n13, A3 => n29, ZN => p(3));
   U44 : MUX2_X1 port map( A => n17, B => n16, S => A(3), Z => n32);
   U45 : MUX2_X1 port map( A => n19, B => n9, S => A(4), Z => n31);
   U46 : NAND3_X1 port map( A1 => n32, A2 => n13, A3 => n31, ZN => p(4));
   U47 : MUX2_X1 port map( A => n17, B => n16, S => A(4), Z => n34);
   U48 : MUX2_X1 port map( A => n20, B => n9, S => A(5), Z => n33);
   U49 : NAND3_X1 port map( A1 => n34, A2 => n13, A3 => n33, ZN => p(5));
   U50 : MUX2_X1 port map( A => n17, B => n16, S => A(5), Z => n36);
   U51 : MUX2_X1 port map( A => n20, B => n9, S => A(6), Z => n35);
   U52 : NAND3_X1 port map( A1 => n36, A2 => n13, A3 => n35, ZN => p(6));
   U53 : MUX2_X1 port map( A => n17, B => n16, S => A(6), Z => n38);
   U54 : MUX2_X1 port map( A => n20, B => n9, S => A(7), Z => n37);
   U55 : NAND3_X1 port map( A1 => n38, A2 => n13, A3 => n37, ZN => p(7));
   U56 : MUX2_X1 port map( A => n21, B => n9, S => A(8), Z => n40);
   U57 : MUX2_X1 port map( A => n17, B => n16, S => A(7), Z => n39);
   U58 : NAND3_X1 port map( A1 => n40, A2 => n12, A3 => n39, ZN => p(8));
   U59 : MUX2_X1 port map( A => n17, B => n16, S => A(8), Z => n42);
   U60 : MUX2_X1 port map( A => n21, B => n9, S => A(9), Z => n41);
   U61 : NAND3_X1 port map( A1 => n42, A2 => n12, A3 => n41, ZN => p(9));
   U62 : MUX2_X1 port map( A => n17, B => n16, S => A(9), Z => n45);
   U63 : NAND2_X1 port map( A1 => n6, A2 => n43, ZN => n76);
   U64 : MUX2_X1 port map( A => n21, B => n89, S => A(10), Z => n44);
   U65 : NAND3_X1 port map( A1 => n45, A2 => n12, A3 => n44, ZN => p(10));
   U66 : MUX2_X1 port map( A => n17, B => n15, S => A(10), Z => n47);
   U67 : MUX2_X1 port map( A => n21, B => n9, S => A(11), Z => n46);
   U68 : NAND3_X1 port map( A1 => n47, A2 => n12, A3 => n46, ZN => p(11));
   U69 : MUX2_X1 port map( A => n17, B => n15, S => A(11), Z => n49);
   U70 : MUX2_X1 port map( A => n19, B => n9, S => A(12), Z => n48);
   U71 : NAND3_X1 port map( A1 => n49, A2 => n12, A3 => n48, ZN => p(12));
   U72 : MUX2_X1 port map( A => n17, B => n15, S => A(12), Z => n51);
   U73 : MUX2_X1 port map( A => n20, B => n9, S => A(13), Z => n50);
   U74 : NAND3_X1 port map( A1 => n51, A2 => n12, A3 => n50, ZN => p(13));
   U75 : MUX2_X1 port map( A => n61, B => n15, S => A(13), Z => n53);
   U76 : MUX2_X1 port map( A => n20, B => n89, S => A(14), Z => n52);
   U77 : NAND3_X1 port map( A1 => n53, A2 => n12, A3 => n52, ZN => p(14));
   U78 : MUX2_X1 port map( A => n61, B => n15, S => A(14), Z => n55);
   U79 : MUX2_X1 port map( A => n19, B => n8, S => A(15), Z => n54);
   U80 : NAND3_X1 port map( A1 => n55, A2 => n12, A3 => n54, ZN => p(15));
   U81 : MUX2_X1 port map( A => n61, B => n15, S => A(15), Z => n57);
   U82 : MUX2_X1 port map( A => n20, B => n76, S => A(16), Z => n56);
   U83 : NAND3_X1 port map( A1 => n57, A2 => n12, A3 => n56, ZN => p(16));
   U84 : MUX2_X1 port map( A => n19, B => n76, S => A(17), Z => n59);
   U85 : MUX2_X1 port map( A => n94, B => n15, S => A(16), Z => n58);
   U86 : NAND3_X1 port map( A1 => n13, A2 => n59, A3 => n58, ZN => p(17));
   U87 : NAND2_X1 port map( A1 => n5, A2 => n60, ZN => n61);
   U88 : MUX2_X1 port map( A => n94, B => n15, S => A(17), Z => n63);
   U89 : MUX2_X1 port map( A => n21, B => n89, S => A(18), Z => n62);
   U90 : NAND3_X1 port map( A1 => n63, A2 => n12, A3 => n62, ZN => p(18));
   U91 : MUX2_X1 port map( A => n17, B => n15, S => A(18), Z => n65);
   U92 : MUX2_X1 port map( A => n20, B => n8, S => A(19), Z => n64);
   U93 : NAND3_X1 port map( A1 => n65, A2 => n12, A3 => n64, ZN => p(19));
   U94 : MUX2_X1 port map( A => n94, B => n15, S => A(19), Z => n67);
   U95 : MUX2_X1 port map( A => n19, B => n89, S => A(20), Z => n66);
   U96 : NAND3_X1 port map( A1 => n67, A2 => n11, A3 => n66, ZN => p(20));
   U97 : MUX2_X1 port map( A => n19, B => n89, S => A(21), Z => n69);
   U98 : MUX2_X1 port map( A => n18, B => n15, S => A(20), Z => n68);
   U99 : NAND3_X1 port map( A1 => n69, A2 => n11, A3 => n68, ZN => p(21));
   U100 : MUX2_X1 port map( A => n18, B => n14, S => A(21), Z => n71);
   U101 : MUX2_X1 port map( A => n19, B => n8, S => A(22), Z => n70);
   U102 : NAND3_X1 port map( A1 => n71, A2 => n11, A3 => n70, ZN => p(22));
   U103 : MUX2_X1 port map( A => n18, B => n14, S => A(22), Z => n73);
   U104 : MUX2_X1 port map( A => n21, B => n8, S => A(23), Z => n72);
   U105 : NAND3_X1 port map( A1 => n73, A2 => n11, A3 => n72, ZN => p(23));
   U106 : MUX2_X1 port map( A => n18, B => n14, S => A(23), Z => n75);
   U107 : MUX2_X1 port map( A => n19, B => n8, S => A(24), Z => n74);
   U108 : NAND3_X1 port map( A1 => n75, A2 => n11, A3 => n74, ZN => p(24));
   U109 : MUX2_X1 port map( A => n61, B => n14, S => A(24), Z => n78);
   U110 : MUX2_X1 port map( A => n21, B => n89, S => A(25), Z => n77);
   U111 : NAND3_X1 port map( A1 => n78, A2 => n11, A3 => n77, ZN => p(25));
   U112 : MUX2_X1 port map( A => n18, B => n14, S => A(25), Z => n80);
   U113 : MUX2_X1 port map( A => n20, B => n8, S => A(26), Z => n79);
   U114 : NAND3_X1 port map( A1 => n80, A2 => n11, A3 => n79, ZN => p(26));
   U115 : MUX2_X1 port map( A => n18, B => n14, S => A(26), Z => n82);
   U116 : MUX2_X1 port map( A => n20, B => n8, S => A(27), Z => n81);
   U117 : NAND3_X1 port map( A1 => n82, A2 => n11, A3 => n81, ZN => p(27));
   U118 : MUX2_X1 port map( A => n18, B => n14, S => A(27), Z => n84);
   U119 : MUX2_X1 port map( A => n21, B => n8, S => A(28), Z => n83);
   U120 : NAND3_X1 port map( A1 => n84, A2 => n11, A3 => n83, ZN => p(28));
   U121 : MUX2_X1 port map( A => n18, B => n14, S => A(28), Z => n86);
   U122 : MUX2_X1 port map( A => n19, B => n8, S => A(29), Z => n85);
   U123 : NAND3_X1 port map( A1 => n86, A2 => n11, A3 => n85, ZN => p(29));
   U124 : MUX2_X1 port map( A => n18, B => n14, S => A(29), Z => n88);
   U125 : MUX2_X1 port map( A => n20, B => n8, S => A(30), Z => n87);
   U126 : NAND3_X1 port map( A1 => n88, A2 => n11, A3 => n87, ZN => p(30));
   U127 : MUX2_X1 port map( A => n18, B => n14, S => A(30), Z => n92);
   U128 : MUX2_X1 port map( A => n21, B => n8, S => A(31), Z => n90);
   U129 : NAND3_X1 port map( A1 => n92, A2 => n12, A3 => n90, ZN => p(31));
   U130 : MUX2_X1 port map( A => n18, B => n14, S => A(31), Z => n95);
   U131 : NAND2_X1 port map( A1 => n21, A2 => n95, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_9 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_9;

architecture SYN_beh of ENC_9 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93 : std_logic;

begin
   
   U3 : BUF_X2 port map( A => n89, Z => n6);
   U4 : BUF_X2 port map( A => n89, Z => n8);
   U5 : BUF_X1 port map( A => n89, Z => n7);
   U6 : OR2_X2 port map( A1 => n19, A2 => b(2), ZN => n87);
   U7 : AND2_X1 port map( A1 => n25, A2 => n26, ZN => n1);
   U8 : BUF_X2 port map( A => n91, Z => n9);
   U9 : BUF_X2 port map( A => n87, Z => n2);
   U10 : BUF_X2 port map( A => n87, Z => n4);
   U11 : CLKBUF_X1 port map( A => n87, Z => n3);
   U12 : NAND3_X1 port map( A1 => n87, A2 => n14, A3 => n1, ZN => n89);
   U13 : BUF_X1 port map( A => n93, Z => n14);
   U14 : CLKBUF_X3 port map( A => n93, Z => n15);
   U15 : BUF_X1 port map( A => n93, Z => n16);
   U16 : BUF_X2 port map( A => n92, Z => n12);
   U17 : BUF_X2 port map( A => n91, Z => n10);
   U18 : BUF_X2 port map( A => n92, Z => n11);
   U19 : CLKBUF_X1 port map( A => n92, Z => n13);
   U20 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n19);
   U21 : CLKBUF_X1 port map( A => n87, Z => n5);
   U22 : INV_X1 port map( A => n18, ZN => n17);
   U23 : INV_X1 port map( A => A(31), ZN => n18);
   U24 : INV_X1 port map( A => b(2), ZN => n22);
   U25 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n21);
   U26 : INV_X1 port map( A => b(0), ZN => n24);
   U27 : INV_X1 port map( A => b(1), ZN => n23);
   U28 : NAND3_X1 port map( A1 => b(2), A2 => n24, A3 => n23, ZN => n92);
   U29 : NAND2_X1 port map( A1 => b(2), A2 => n21, ZN => n25);
   U30 : MUX2_X1 port map( A => n25, B => n2, S => A(0), Z => n20);
   U31 : OAI211_X1 port map( C1 => n22, C2 => n21, A => n11, B => n20, ZN => 
                           p(0));
   U32 : NAND3_X1 port map( A1 => b(1), A2 => n22, A3 => b(0), ZN => n93);
   U33 : MUX2_X1 port map( A => n11, B => n16, S => A(0), Z => n28);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n23, ZN => n26);
   U35 : NAND2_X1 port map( A1 => b(2), A2 => n26, ZN => n91);
   U36 : MUX2_X1 port map( A => n10, B => n2, S => A(1), Z => n27);
   U37 : NAND3_X1 port map( A1 => n28, A2 => n8, A3 => n27, ZN => p(1));
   U38 : MUX2_X1 port map( A => n11, B => n15, S => A(1), Z => n30);
   U39 : MUX2_X1 port map( A => n10, B => n5, S => A(2), Z => n29);
   U40 : NAND3_X1 port map( A1 => n30, A2 => n6, A3 => n29, ZN => p(2));
   U41 : MUX2_X1 port map( A => n11, B => n16, S => A(2), Z => n32);
   U42 : MUX2_X1 port map( A => n10, B => n2, S => A(3), Z => n31);
   U43 : NAND3_X1 port map( A1 => n32, A2 => n8, A3 => n31, ZN => p(3));
   U44 : MUX2_X1 port map( A => n11, B => n16, S => A(3), Z => n34);
   U45 : MUX2_X1 port map( A => n10, B => n4, S => A(4), Z => n33);
   U46 : NAND3_X1 port map( A1 => n34, A2 => n6, A3 => n33, ZN => p(4));
   U47 : MUX2_X1 port map( A => n11, B => n15, S => A(4), Z => n36);
   U48 : MUX2_X1 port map( A => n10, B => n4, S => A(5), Z => n35);
   U49 : NAND3_X1 port map( A1 => n36, A2 => n8, A3 => n35, ZN => p(5));
   U50 : MUX2_X1 port map( A => n11, B => n16, S => A(5), Z => n38);
   U51 : MUX2_X1 port map( A => n10, B => n2, S => A(6), Z => n37);
   U52 : NAND3_X1 port map( A1 => n38, A2 => n6, A3 => n37, ZN => p(6));
   U53 : MUX2_X1 port map( A => n11, B => n15, S => A(6), Z => n40);
   U54 : MUX2_X1 port map( A => n10, B => n2, S => A(7), Z => n39);
   U55 : NAND3_X1 port map( A1 => n40, A2 => n6, A3 => n39, ZN => p(7));
   U56 : MUX2_X1 port map( A => n12, B => n15, S => A(7), Z => n42);
   U57 : MUX2_X1 port map( A => n10, B => n5, S => A(8), Z => n41);
   U58 : NAND3_X1 port map( A1 => n42, A2 => n8, A3 => n41, ZN => p(8));
   U59 : MUX2_X1 port map( A => n11, B => n15, S => A(8), Z => n44);
   U60 : MUX2_X1 port map( A => n10, B => n4, S => A(9), Z => n43);
   U61 : NAND3_X1 port map( A1 => n44, A2 => n6, A3 => n43, ZN => p(9));
   U62 : MUX2_X1 port map( A => n10, B => n4, S => A(10), Z => n46);
   U63 : MUX2_X1 port map( A => n11, B => n15, S => A(9), Z => n45);
   U64 : NAND3_X1 port map( A1 => n46, A2 => n7, A3 => n45, ZN => p(10));
   U65 : MUX2_X1 port map( A => n11, B => n16, S => A(10), Z => n48);
   U66 : MUX2_X1 port map( A => n10, B => n2, S => A(11), Z => n47);
   U67 : NAND3_X1 port map( A1 => n48, A2 => n8, A3 => n47, ZN => p(11));
   U68 : MUX2_X1 port map( A => n11, B => n16, S => A(11), Z => n50);
   U69 : MUX2_X1 port map( A => n10, B => n4, S => A(12), Z => n49);
   U70 : NAND3_X1 port map( A1 => n50, A2 => n8, A3 => n49, ZN => p(12));
   U71 : MUX2_X1 port map( A => n10, B => n5, S => A(13), Z => n52);
   U72 : MUX2_X1 port map( A => n11, B => n15, S => A(12), Z => n51);
   U73 : NAND3_X1 port map( A1 => n52, A2 => n7, A3 => n51, ZN => p(13));
   U74 : MUX2_X1 port map( A => n10, B => n3, S => A(14), Z => n54);
   U75 : MUX2_X1 port map( A => n12, B => n16, S => A(13), Z => n53);
   U76 : NAND3_X1 port map( A1 => n7, A2 => n54, A3 => n53, ZN => p(14));
   U77 : MUX2_X1 port map( A => n10, B => n4, S => A(15), Z => n56);
   U78 : MUX2_X1 port map( A => n12, B => n15, S => A(14), Z => n55);
   U79 : NAND3_X1 port map( A1 => n56, A2 => n6, A3 => n55, ZN => p(15));
   U80 : MUX2_X1 port map( A => n12, B => n16, S => A(15), Z => n58);
   U81 : MUX2_X1 port map( A => n10, B => n2, S => A(16), Z => n57);
   U82 : NAND3_X1 port map( A1 => n58, A2 => n6, A3 => n57, ZN => p(16));
   U83 : MUX2_X1 port map( A => n12, B => n15, S => A(16), Z => n60);
   U84 : MUX2_X1 port map( A => n9, B => n2, S => A(17), Z => n59);
   U85 : NAND3_X1 port map( A1 => n60, A2 => n6, A3 => n59, ZN => p(17));
   U86 : MUX2_X1 port map( A => n12, B => n15, S => A(17), Z => n62);
   U87 : MUX2_X1 port map( A => n9, B => n2, S => A(18), Z => n61);
   U88 : NAND3_X1 port map( A1 => n62, A2 => n7, A3 => n61, ZN => p(18));
   U89 : MUX2_X1 port map( A => n9, B => n4, S => A(19), Z => n64);
   U90 : MUX2_X1 port map( A => n12, B => n15, S => A(18), Z => n63);
   U91 : NAND3_X1 port map( A1 => n64, A2 => n63, A3 => n6, ZN => p(19));
   U92 : MUX2_X1 port map( A => n12, B => n15, S => A(19), Z => n66);
   U93 : MUX2_X1 port map( A => n9, B => n4, S => A(20), Z => n65);
   U94 : NAND3_X1 port map( A1 => n66, A2 => n8, A3 => n65, ZN => p(20));
   U95 : MUX2_X1 port map( A => n12, B => n16, S => A(20), Z => n68);
   U96 : MUX2_X1 port map( A => n9, B => n4, S => A(21), Z => n67);
   U97 : NAND3_X1 port map( A1 => n68, A2 => n8, A3 => n67, ZN => p(21));
   U98 : MUX2_X1 port map( A => n9, B => n2, S => A(22), Z => n70);
   U99 : MUX2_X1 port map( A => n12, B => n16, S => A(21), Z => n69);
   U100 : NAND3_X1 port map( A1 => n70, A2 => n7, A3 => n69, ZN => p(22));
   U101 : MUX2_X1 port map( A => n12, B => n16, S => A(22), Z => n72);
   U102 : MUX2_X1 port map( A => n9, B => n4, S => A(23), Z => n71);
   U103 : NAND3_X1 port map( A1 => n72, A2 => n8, A3 => n71, ZN => p(23));
   U104 : MUX2_X1 port map( A => n12, B => n16, S => A(23), Z => n74);
   U105 : MUX2_X1 port map( A => n9, B => n4, S => A(24), Z => n73);
   U106 : NAND3_X1 port map( A1 => n74, A2 => n6, A3 => n73, ZN => p(24));
   U107 : MUX2_X1 port map( A => n12, B => n15, S => A(24), Z => n76);
   U108 : MUX2_X1 port map( A => n9, B => n5, S => A(25), Z => n75);
   U109 : NAND3_X1 port map( A1 => n76, A2 => n6, A3 => n75, ZN => p(25));
   U110 : MUX2_X1 port map( A => n12, B => n15, S => A(25), Z => n78);
   U111 : MUX2_X1 port map( A => n9, B => n4, S => A(26), Z => n77);
   U112 : NAND3_X1 port map( A1 => n78, A2 => n8, A3 => n77, ZN => p(26));
   U113 : MUX2_X1 port map( A => n12, B => n16, S => A(26), Z => n80);
   U114 : MUX2_X1 port map( A => n9, B => n2, S => A(27), Z => n79);
   U115 : NAND3_X1 port map( A1 => n80, A2 => n8, A3 => n79, ZN => p(27));
   U116 : MUX2_X1 port map( A => n12, B => n15, S => A(27), Z => n82);
   U117 : MUX2_X1 port map( A => n9, B => n5, S => A(28), Z => n81);
   U118 : NAND3_X1 port map( A1 => n82, A2 => n8, A3 => n81, ZN => p(28));
   U119 : MUX2_X1 port map( A => n13, B => n15, S => A(28), Z => n84);
   U120 : MUX2_X1 port map( A => n9, B => n2, S => A(29), Z => n83);
   U121 : NAND3_X1 port map( A1 => n84, A2 => n6, A3 => n83, ZN => p(29));
   U122 : MUX2_X1 port map( A => n13, B => n16, S => A(29), Z => n86);
   U123 : MUX2_X1 port map( A => n9, B => n2, S => A(30), Z => n85);
   U124 : NAND3_X1 port map( A1 => n86, A2 => n6, A3 => n85, ZN => p(30));
   U125 : MUX2_X1 port map( A => n11, B => n15, S => A(30), Z => n90);
   U126 : MUX2_X1 port map( A => n9, B => n4, S => n17, Z => n88);
   U127 : NAND3_X1 port map( A1 => n90, A2 => n6, A3 => n88, ZN => p(31));
   U128 : OAI221_X1 port map( B1 => n18, B2 => n15, C1 => n17, C2 => n11, A => 
                           n9, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_8 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_8;

architecture SYN_beh of ENC_8 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90 : std_logic;

begin
   
   U3 : BUF_X2 port map( A => n84, Z => n4);
   U4 : BUF_X1 port map( A => n84, Z => n2);
   U5 : OR2_X2 port map( A1 => n19, A2 => b(2), ZN => n84);
   U6 : CLKBUF_X1 port map( A => b(0), Z => n1);
   U7 : BUF_X2 port map( A => n84, Z => n3);
   U8 : BUF_X1 port map( A => n88, Z => n8);
   U9 : BUF_X1 port map( A => n86, Z => n5);
   U10 : BUF_X1 port map( A => n86, Z => n6);
   U11 : BUF_X2 port map( A => n88, Z => n9);
   U12 : BUF_X2 port map( A => n89, Z => n11);
   U13 : BUF_X2 port map( A => n90, Z => n14);
   U14 : BUF_X2 port map( A => n89, Z => n10);
   U15 : BUF_X1 port map( A => n90, Z => n13);
   U16 : BUF_X1 port map( A => n86, Z => n7);
   U17 : MUX2_X1 port map( A => n12, B => n13, S => A(29), Z => n83);
   U18 : MUX2_X1 port map( A => n12, B => n13, S => A(30), Z => n87);
   U19 : CLKBUF_X1 port map( A => n89, Z => n12);
   U20 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n19);
   U21 : INV_X1 port map( A => n16, ZN => n15);
   U22 : INV_X1 port map( A => A(31), ZN => n16);
   U23 : INV_X1 port map( A => b(2), ZN => n22);
   U24 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n21);
   U25 : INV_X1 port map( A => b(0), ZN => n18);
   U26 : INV_X1 port map( A => b(1), ZN => n17);
   U27 : NAND3_X1 port map( A1 => b(2), A2 => n18, A3 => n17, ZN => n89);
   U28 : NAND2_X1 port map( A1 => b(2), A2 => n21, ZN => n23);
   U29 : MUX2_X1 port map( A => n23, B => n4, S => A(0), Z => n20);
   U30 : OAI211_X1 port map( C1 => n22, C2 => n21, A => n10, B => n20, ZN => 
                           p(0));
   U31 : NAND2_X1 port map( A1 => b(1), A2 => n1, ZN => n90);
   U32 : MUX2_X1 port map( A => n10, B => n13, S => A(0), Z => n25);
   U33 : NAND2_X1 port map( A1 => b(2), A2 => n23, ZN => n86);
   U34 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => b(2), ZN => n88);
   U35 : MUX2_X1 port map( A => n9, B => n4, S => A(1), Z => n24);
   U36 : NAND3_X1 port map( A1 => n25, A2 => n5, A3 => n24, ZN => p(1));
   U37 : MUX2_X1 port map( A => n10, B => n13, S => A(1), Z => n27);
   U38 : MUX2_X1 port map( A => n9, B => n2, S => A(2), Z => n26);
   U39 : NAND3_X1 port map( A1 => n27, A2 => n7, A3 => n26, ZN => p(2));
   U40 : MUX2_X1 port map( A => n10, B => n13, S => A(2), Z => n29);
   U41 : MUX2_X1 port map( A => n9, B => n4, S => A(3), Z => n28);
   U42 : NAND3_X1 port map( A1 => n29, A2 => n7, A3 => n28, ZN => p(3));
   U43 : MUX2_X1 port map( A => n10, B => n13, S => A(3), Z => n31);
   U44 : MUX2_X1 port map( A => n9, B => n2, S => A(4), Z => n30);
   U45 : NAND3_X1 port map( A1 => n31, A2 => n7, A3 => n30, ZN => p(4));
   U46 : MUX2_X1 port map( A => n10, B => n13, S => A(4), Z => n33);
   U47 : MUX2_X1 port map( A => n9, B => n2, S => A(5), Z => n32);
   U48 : NAND3_X1 port map( A1 => n33, A2 => n7, A3 => n32, ZN => p(5));
   U49 : MUX2_X1 port map( A => n10, B => n13, S => A(5), Z => n35);
   U50 : MUX2_X1 port map( A => n9, B => n4, S => A(6), Z => n34);
   U51 : NAND3_X1 port map( A1 => n35, A2 => n7, A3 => n34, ZN => p(6));
   U52 : MUX2_X1 port map( A => n9, B => n3, S => A(7), Z => n37);
   U53 : MUX2_X1 port map( A => n10, B => n14, S => A(6), Z => n36);
   U54 : NAND3_X1 port map( A1 => n37, A2 => n7, A3 => n36, ZN => p(7));
   U55 : MUX2_X1 port map( A => n9, B => n2, S => A(8), Z => n39);
   U56 : MUX2_X1 port map( A => n11, B => n13, S => A(7), Z => n38);
   U57 : NAND3_X1 port map( A1 => n39, A2 => n6, A3 => n38, ZN => p(8));
   U58 : MUX2_X1 port map( A => n10, B => n13, S => A(8), Z => n41);
   U59 : MUX2_X1 port map( A => n9, B => n4, S => A(9), Z => n40);
   U60 : NAND3_X1 port map( A1 => n41, A2 => n6, A3 => n40, ZN => p(9));
   U61 : MUX2_X1 port map( A => n9, B => n3, S => A(10), Z => n43);
   U62 : MUX2_X1 port map( A => n10, B => n14, S => A(9), Z => n42);
   U63 : NAND3_X1 port map( A1 => n7, A2 => n43, A3 => n42, ZN => p(10));
   U64 : MUX2_X1 port map( A => n10, B => n13, S => A(10), Z => n45);
   U65 : MUX2_X1 port map( A => n9, B => n4, S => A(11), Z => n44);
   U66 : NAND3_X1 port map( A1 => n45, A2 => n6, A3 => n44, ZN => p(11));
   U67 : MUX2_X1 port map( A => n10, B => n14, S => A(11), Z => n47);
   U68 : MUX2_X1 port map( A => n9, B => n2, S => A(12), Z => n46);
   U69 : NAND3_X1 port map( A1 => n47, A2 => n6, A3 => n46, ZN => p(12));
   U70 : MUX2_X1 port map( A => n9, B => n2, S => A(13), Z => n49);
   U71 : MUX2_X1 port map( A => n10, B => n14, S => A(12), Z => n48);
   U72 : NAND3_X1 port map( A1 => n49, A2 => n6, A3 => n48, ZN => p(13));
   U73 : MUX2_X1 port map( A => n9, B => n3, S => A(14), Z => n51);
   U74 : MUX2_X1 port map( A => n10, B => n14, S => A(13), Z => n50);
   U75 : NAND3_X1 port map( A1 => n51, A2 => n50, A3 => n5, ZN => p(14));
   U76 : MUX2_X1 port map( A => n11, B => n14, S => A(14), Z => n53);
   U77 : MUX2_X1 port map( A => n9, B => n3, S => A(15), Z => n52);
   U78 : NAND3_X1 port map( A1 => n52, A2 => n53, A3 => n5, ZN => p(15));
   U79 : MUX2_X1 port map( A => n9, B => n3, S => A(16), Z => n55);
   U80 : MUX2_X1 port map( A => n11, B => n14, S => A(15), Z => n54);
   U81 : NAND3_X1 port map( A1 => n55, A2 => n6, A3 => n54, ZN => p(16));
   U82 : MUX2_X1 port map( A => n11, B => n13, S => A(16), Z => n57);
   U83 : MUX2_X1 port map( A => n8, B => n4, S => A(17), Z => n56);
   U84 : NAND3_X1 port map( A1 => n57, A2 => n6, A3 => n56, ZN => p(17));
   U85 : MUX2_X1 port map( A => n11, B => n13, S => A(17), Z => n59);
   U86 : MUX2_X1 port map( A => n8, B => n4, S => A(18), Z => n58);
   U87 : NAND3_X1 port map( A1 => n59, A2 => n6, A3 => n58, ZN => p(18));
   U88 : MUX2_X1 port map( A => n11, B => n14, S => A(18), Z => n61);
   U89 : MUX2_X1 port map( A => n8, B => n2, S => A(19), Z => n60);
   U90 : NAND3_X1 port map( A1 => n61, A2 => n6, A3 => n60, ZN => p(19));
   U91 : MUX2_X1 port map( A => n11, B => n14, S => A(19), Z => n63);
   U92 : MUX2_X1 port map( A => n8, B => n3, S => A(20), Z => n62);
   U93 : NAND3_X1 port map( A1 => n63, A2 => n6, A3 => n62, ZN => p(20));
   U94 : MUX2_X1 port map( A => n11, B => n13, S => A(20), Z => n65);
   U95 : MUX2_X1 port map( A => n8, B => n4, S => A(21), Z => n64);
   U96 : NAND3_X1 port map( A1 => n65, A2 => n5, A3 => n64, ZN => p(21));
   U97 : MUX2_X1 port map( A => n11, B => n13, S => A(21), Z => n67);
   U98 : MUX2_X1 port map( A => n8, B => n4, S => A(22), Z => n66);
   U99 : NAND3_X1 port map( A1 => n67, A2 => n6, A3 => n66, ZN => p(22));
   U100 : MUX2_X1 port map( A => n11, B => n13, S => A(22), Z => n69);
   U101 : MUX2_X1 port map( A => n8, B => n4, S => A(23), Z => n68);
   U102 : NAND3_X1 port map( A1 => n69, A2 => n5, A3 => n68, ZN => p(23));
   U103 : MUX2_X1 port map( A => n11, B => n13, S => A(23), Z => n71);
   U104 : MUX2_X1 port map( A => n8, B => n2, S => A(24), Z => n70);
   U105 : NAND3_X1 port map( A1 => n71, A2 => n5, A3 => n70, ZN => p(24));
   U106 : MUX2_X1 port map( A => n11, B => n13, S => A(24), Z => n73);
   U107 : MUX2_X1 port map( A => n8, B => n4, S => A(25), Z => n72);
   U108 : NAND3_X1 port map( A1 => n73, A2 => n5, A3 => n72, ZN => p(25));
   U109 : MUX2_X1 port map( A => n11, B => n13, S => A(25), Z => n75);
   U110 : MUX2_X1 port map( A => n8, B => n2, S => A(26), Z => n74);
   U111 : NAND3_X1 port map( A1 => n75, A2 => n5, A3 => n74, ZN => p(26));
   U112 : MUX2_X1 port map( A => n11, B => n13, S => A(26), Z => n77);
   U113 : MUX2_X1 port map( A => n8, B => n2, S => A(27), Z => n76);
   U114 : NAND3_X1 port map( A1 => n77, A2 => n5, A3 => n76, ZN => p(27));
   U115 : MUX2_X1 port map( A => n11, B => n13, S => A(27), Z => n79);
   U116 : MUX2_X1 port map( A => n8, B => n4, S => A(28), Z => n78);
   U117 : NAND3_X1 port map( A1 => n79, A2 => n5, A3 => n78, ZN => p(28));
   U118 : MUX2_X1 port map( A => n11, B => n13, S => A(28), Z => n81);
   U119 : MUX2_X1 port map( A => n8, B => n4, S => A(29), Z => n80);
   U120 : NAND3_X1 port map( A1 => n81, A2 => n5, A3 => n80, ZN => p(29));
   U121 : MUX2_X1 port map( A => n8, B => n2, S => A(30), Z => n82);
   U122 : NAND3_X1 port map( A1 => n83, A2 => n5, A3 => n82, ZN => p(30));
   U123 : MUX2_X1 port map( A => n8, B => n4, S => n15, Z => n85);
   U124 : NAND3_X1 port map( A1 => n87, A2 => n6, A3 => n85, ZN => p(31));
   U125 : OAI221_X1 port map( B1 => n16, B2 => n13, C1 => n15, C2 => n10, A => 
                           n8, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_7 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_7;

architecture SYN_beh of ENC_7 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91 : std_logic;

begin
   
   U3 : NAND3_X1 port map( A1 => n56, A2 => n7, A3 => n55, ZN => p(16));
   U4 : OR2_X1 port map( A1 => n20, A2 => b(2), ZN => n1);
   U5 : OR2_X1 port map( A1 => n20, A2 => b(2), ZN => n85);
   U6 : BUF_X1 port map( A => n85, Z => n4);
   U7 : BUF_X1 port map( A => n85, Z => n5);
   U8 : BUF_X2 port map( A => n90, Z => n12);
   U9 : CLKBUF_X1 port map( A => b(0), Z => n2);
   U10 : BUF_X2 port map( A => n85, Z => n3);
   U11 : BUF_X1 port map( A => n89, Z => n9);
   U12 : BUF_X1 port map( A => n87, Z => n6);
   U13 : BUF_X1 port map( A => n87, Z => n7);
   U14 : BUF_X2 port map( A => n89, Z => n10);
   U15 : BUF_X2 port map( A => n91, Z => n15);
   U16 : BUF_X2 port map( A => n90, Z => n11);
   U17 : BUF_X1 port map( A => n91, Z => n14);
   U18 : BUF_X1 port map( A => n87, Z => n8);
   U19 : MUX2_X1 port map( A => n12, B => n14, S => A(28), Z => n82);
   U20 : MUX2_X1 port map( A => n13, B => n14, S => A(29), Z => n84);
   U21 : MUX2_X1 port map( A => n13, B => n14, S => A(30), Z => n88);
   U22 : MUX2_X1 port map( A => n12, B => n14, S => A(27), Z => n80);
   U23 : CLKBUF_X1 port map( A => n90, Z => n13);
   U24 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n20);
   U25 : INV_X1 port map( A => n17, ZN => n16);
   U26 : INV_X1 port map( A => A(31), ZN => n17);
   U27 : INV_X1 port map( A => b(2), ZN => n23);
   U28 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n22);
   U29 : INV_X1 port map( A => b(0), ZN => n19);
   U30 : INV_X1 port map( A => b(1), ZN => n18);
   U31 : NAND3_X1 port map( A1 => b(2), A2 => n19, A3 => n18, ZN => n90);
   U32 : NAND2_X1 port map( A1 => b(2), A2 => n22, ZN => n24);
   U33 : MUX2_X1 port map( A => n24, B => n1, S => A(0), Z => n21);
   U34 : OAI211_X1 port map( C1 => n23, C2 => n22, A => n11, B => n21, ZN => 
                           p(0));
   U35 : NAND2_X1 port map( A1 => b(1), A2 => n2, ZN => n91);
   U36 : MUX2_X1 port map( A => n11, B => n14, S => A(0), Z => n26);
   U37 : NAND2_X1 port map( A1 => b(2), A2 => n24, ZN => n87);
   U38 : OAI21_X1 port map( B1 => b(0), B2 => b(1), A => b(2), ZN => n89);
   U39 : MUX2_X1 port map( A => n10, B => n3, S => A(1), Z => n25);
   U40 : NAND3_X1 port map( A1 => n26, A2 => n6, A3 => n25, ZN => p(1));
   U41 : MUX2_X1 port map( A => n11, B => n15, S => A(1), Z => n28);
   U42 : MUX2_X1 port map( A => n10, B => n3, S => A(2), Z => n27);
   U43 : NAND3_X1 port map( A1 => n28, A2 => n8, A3 => n27, ZN => p(2));
   U44 : MUX2_X1 port map( A => n11, B => n15, S => A(2), Z => n30);
   U45 : MUX2_X1 port map( A => n10, B => n4, S => A(3), Z => n29);
   U46 : NAND3_X1 port map( A1 => n30, A2 => n8, A3 => n29, ZN => p(3));
   U47 : MUX2_X1 port map( A => n11, B => n15, S => A(3), Z => n32);
   U48 : MUX2_X1 port map( A => n10, B => n85, S => A(4), Z => n31);
   U49 : NAND3_X1 port map( A1 => n32, A2 => n8, A3 => n31, ZN => p(4));
   U50 : MUX2_X1 port map( A => n10, B => n5, S => A(5), Z => n34);
   U51 : MUX2_X1 port map( A => n11, B => n15, S => A(4), Z => n33);
   U52 : NAND3_X1 port map( A1 => n34, A2 => n8, A3 => n33, ZN => p(5));
   U53 : MUX2_X1 port map( A => n11, B => n15, S => A(5), Z => n36);
   U54 : MUX2_X1 port map( A => n10, B => n1, S => A(6), Z => n35);
   U55 : NAND3_X1 port map( A1 => n36, A2 => n8, A3 => n35, ZN => p(6));
   U56 : MUX2_X1 port map( A => n11, B => n15, S => A(6), Z => n38);
   U57 : MUX2_X1 port map( A => n10, B => n4, S => A(7), Z => n37);
   U58 : NAND3_X1 port map( A1 => n38, A2 => n8, A3 => n37, ZN => p(7));
   U59 : MUX2_X1 port map( A => n10, B => n85, S => A(8), Z => n40);
   U60 : MUX2_X1 port map( A => n12, B => n15, S => A(7), Z => n39);
   U61 : NAND3_X1 port map( A1 => n8, A2 => n40, A3 => n39, ZN => p(8));
   U62 : MUX2_X1 port map( A => n11, B => n15, S => A(8), Z => n42);
   U63 : MUX2_X1 port map( A => n10, B => n1, S => A(9), Z => n41);
   U64 : NAND3_X1 port map( A1 => n42, A2 => n7, A3 => n41, ZN => p(9));
   U65 : MUX2_X1 port map( A => n11, B => n15, S => A(9), Z => n44);
   U66 : MUX2_X1 port map( A => n10, B => n85, S => A(10), Z => n43);
   U67 : NAND3_X1 port map( A1 => n44, A2 => n7, A3 => n43, ZN => p(10));
   U68 : MUX2_X1 port map( A => n10, B => n1, S => A(11), Z => n46);
   U69 : MUX2_X1 port map( A => n11, B => n15, S => A(10), Z => n45);
   U70 : NAND3_X1 port map( A1 => n46, A2 => n45, A3 => n6, ZN => p(11));
   U71 : MUX2_X1 port map( A => n10, B => n1, S => A(12), Z => n48);
   U72 : MUX2_X1 port map( A => n11, B => n15, S => A(11), Z => n47);
   U73 : NAND3_X1 port map( A1 => n48, A2 => n47, A3 => n6, ZN => p(12));
   U74 : MUX2_X1 port map( A => n11, B => n15, S => A(12), Z => n50);
   U75 : MUX2_X1 port map( A => n10, B => n1, S => A(13), Z => n49);
   U76 : NAND3_X1 port map( A1 => n50, A2 => n7, A3 => n49, ZN => p(13));
   U77 : MUX2_X1 port map( A => n11, B => n15, S => A(13), Z => n52);
   U78 : MUX2_X1 port map( A => n10, B => n85, S => A(14), Z => n51);
   U79 : NAND3_X1 port map( A1 => n52, A2 => n7, A3 => n51, ZN => p(14));
   U80 : MUX2_X1 port map( A => n12, B => n15, S => A(14), Z => n54);
   U81 : MUX2_X1 port map( A => n10, B => n1, S => A(15), Z => n53);
   U82 : NAND3_X1 port map( A1 => n54, A2 => n7, A3 => n53, ZN => p(15));
   U83 : MUX2_X1 port map( A => n12, B => n15, S => A(15), Z => n56);
   U84 : MUX2_X1 port map( A => n10, B => n85, S => A(16), Z => n55);
   U85 : MUX2_X1 port map( A => n12, B => n15, S => A(16), Z => n58);
   U86 : MUX2_X1 port map( A => n9, B => n85, S => A(17), Z => n57);
   U87 : NAND3_X1 port map( A1 => n58, A2 => n7, A3 => n57, ZN => p(17));
   U88 : MUX2_X1 port map( A => n12, B => n14, S => A(17), Z => n60);
   U89 : MUX2_X1 port map( A => n9, B => n85, S => A(18), Z => n59);
   U90 : NAND3_X1 port map( A1 => n60, A2 => n7, A3 => n59, ZN => p(18));
   U91 : MUX2_X1 port map( A => n12, B => n14, S => A(18), Z => n62);
   U92 : MUX2_X1 port map( A => n9, B => n5, S => A(19), Z => n61);
   U93 : NAND3_X1 port map( A1 => n62, A2 => n7, A3 => n61, ZN => p(19));
   U94 : MUX2_X1 port map( A => n12, B => n14, S => A(19), Z => n64);
   U95 : MUX2_X1 port map( A => n9, B => n1, S => A(20), Z => n63);
   U96 : NAND3_X1 port map( A1 => n64, A2 => n7, A3 => n63, ZN => p(20));
   U97 : MUX2_X1 port map( A => n12, B => n14, S => A(20), Z => n66);
   U98 : MUX2_X1 port map( A => n9, B => n85, S => A(21), Z => n65);
   U99 : NAND3_X1 port map( A1 => n66, A2 => n7, A3 => n65, ZN => p(21));
   U100 : MUX2_X1 port map( A => n12, B => n14, S => A(21), Z => n68);
   U101 : MUX2_X1 port map( A => n9, B => n85, S => A(22), Z => n67);
   U102 : NAND3_X1 port map( A1 => n68, A2 => n6, A3 => n67, ZN => p(22));
   U103 : MUX2_X1 port map( A => n12, B => n14, S => A(22), Z => n70);
   U104 : MUX2_X1 port map( A => n9, B => n4, S => A(23), Z => n69);
   U105 : NAND3_X1 port map( A1 => n70, A2 => n6, A3 => n69, ZN => p(23));
   U106 : MUX2_X1 port map( A => n12, B => n14, S => A(23), Z => n72);
   U107 : MUX2_X1 port map( A => n9, B => n3, S => A(24), Z => n71);
   U108 : NAND3_X1 port map( A1 => n72, A2 => n6, A3 => n71, ZN => p(24));
   U109 : MUX2_X1 port map( A => n12, B => n14, S => A(24), Z => n74);
   U110 : MUX2_X1 port map( A => n9, B => n3, S => A(25), Z => n73);
   U111 : NAND3_X1 port map( A1 => n74, A2 => n6, A3 => n73, ZN => p(25));
   U112 : MUX2_X1 port map( A => n12, B => n14, S => A(25), Z => n76);
   U113 : MUX2_X1 port map( A => n9, B => n3, S => A(26), Z => n75);
   U114 : NAND3_X1 port map( A1 => n76, A2 => n6, A3 => n75, ZN => p(26));
   U115 : MUX2_X1 port map( A => n12, B => n14, S => A(26), Z => n78);
   U116 : MUX2_X1 port map( A => n9, B => n3, S => A(27), Z => n77);
   U117 : NAND3_X1 port map( A1 => n78, A2 => n6, A3 => n77, ZN => p(27));
   U118 : MUX2_X1 port map( A => n9, B => n3, S => A(28), Z => n79);
   U119 : NAND3_X1 port map( A1 => n80, A2 => n6, A3 => n79, ZN => p(28));
   U120 : MUX2_X1 port map( A => n9, B => n3, S => A(29), Z => n81);
   U121 : NAND3_X1 port map( A1 => n82, A2 => n6, A3 => n81, ZN => p(29));
   U122 : MUX2_X1 port map( A => n9, B => n3, S => A(30), Z => n83);
   U123 : NAND3_X1 port map( A1 => n84, A2 => n6, A3 => n83, ZN => p(30));
   U124 : MUX2_X1 port map( A => n9, B => n3, S => n16, Z => n86);
   U125 : NAND3_X1 port map( A1 => n88, A2 => n7, A3 => n86, ZN => p(31));
   U126 : OAI221_X1 port map( B1 => n17, B2 => n14, C1 => n16, C2 => n11, A => 
                           n9, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_6 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_6;

architecture SYN_beh of ENC_6 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29488, net29492, net29502, net29521, net29523, net31021, net31019,
      net31029, net31027, net31025, net31033, net31031, net31039, net31037, 
      net31035, net31045, net29526, net29525, net29490, net29455, net29452, 
      net29451, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   U3 : CLKBUF_X1 port map( A => net29452, Z => net31025);
   U4 : BUF_X2 port map( A => net29452, Z => net31027);
   U5 : OR2_X2 port map( A1 => b(2), A2 => n4, ZN => n2);
   U6 : BUF_X2 port map( A => net29455, Z => net31037);
   U7 : OR2_X1 port map( A1 => b(2), A2 => n4, ZN => n1);
   U8 : OR2_X2 port map( A1 => b(2), A2 => n4, ZN => net31045);
   U9 : NAND3_X1 port map( A1 => n5, A2 => net31037, A3 => net29490, ZN => 
                           p(14));
   U10 : MUX2_X1 port map( A => net31027, B => net31021, S => A(14), Z => 
                           net29488);
   U11 : MUX2_X1 port map( A => net31031, B => n2, S => A(14), Z => n5);
   U12 : XNOR2_X1 port map( A => b(1), B => b(0), ZN => n4);
   U13 : OR2_X1 port map( A1 => b(1), A2 => b(0), ZN => n6);
   U14 : NAND2_X1 port map( A1 => n6, A2 => b(2), ZN => n3);
   U15 : CLKBUF_X1 port map( A => n3, Z => n7);
   U16 : BUF_X2 port map( A => n3, Z => net31031);
   U17 : BUF_X1 port map( A => n3, Z => net31033);
   U18 : MUX2_X1 port map( A => net31025, B => net31021, S => A(13), Z => 
                           net29490);
   U19 : BUF_X2 port map( A => net29451, Z => net31021);
   U20 : NAND2_X1 port map( A1 => b(2), A2 => net29521, ZN => net29455);
   U21 : BUF_X1 port map( A => net29455, Z => net31039);
   U22 : BUF_X1 port map( A => net29455, Z => net31035);
   U23 : MUX2_X1 port map( A => net31033, B => n1, S => A(13), Z => net29492);
   U24 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => net29451);
   U25 : BUF_X1 port map( A => net29451, Z => net31019);
   U26 : NAND3_X1 port map( A1 => b(2), A2 => net29525, A3 => net29526, ZN => 
                           net29452);
   U27 : CLKBUF_X1 port map( A => net29452, Z => net31029);
   U28 : INV_X1 port map( A => b(1), ZN => net29526);
   U29 : INV_X1 port map( A => b(0), ZN => net29525);
   U30 : MUX2_X1 port map( A => net29521, B => net31045, S => A(0), Z => 
                           net29523);
   U31 : MUX2_X1 port map( A => net31027, B => net31019, S => A(26), Z => n62);
   U32 : MUX2_X1 port map( A => net31027, B => net31019, S => A(27), Z => n64);
   U33 : MUX2_X1 port map( A => net31027, B => net31019, S => A(28), Z => n66);
   U34 : MUX2_X1 port map( A => net31027, B => net31019, S => A(29), Z => n68);
   U35 : MUX2_X1 port map( A => net31027, B => net31019, S => A(30), Z => n70);
   U36 : MUX2_X1 port map( A => net31027, B => net31019, S => A(25), Z => n60);
   U37 : INV_X1 port map( A => n9, ZN => n8);
   U38 : INV_X1 port map( A => A(31), ZN => n9);
   U39 : INV_X1 port map( A => b(2), ZN => net29502);
   U40 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n10);
   U41 : NAND2_X1 port map( A1 => b(2), A2 => n10, ZN => net29521);
   U42 : OAI211_X1 port map( C1 => net29502, C2 => n10, A => net31029, B => 
                           net29523, ZN => p(0));
   U43 : MUX2_X1 port map( A => net31029, B => net31019, S => A(0), Z => n12);
   U44 : MUX2_X1 port map( A => net31031, B => n1, S => A(1), Z => n11);
   U45 : NAND3_X1 port map( A1 => n12, A2 => net31035, A3 => n11, ZN => p(1));
   U46 : MUX2_X1 port map( A => net31027, B => net31021, S => A(1), Z => n14);
   U47 : MUX2_X1 port map( A => net31033, B => net31045, S => A(2), Z => n13);
   U48 : NAND3_X1 port map( A1 => n14, A2 => net31039, A3 => n13, ZN => p(2));
   U49 : MUX2_X1 port map( A => net31025, B => net31021, S => A(2), Z => n16);
   U50 : MUX2_X1 port map( A => net31033, B => net31045, S => A(3), Z => n15);
   U51 : NAND3_X1 port map( A1 => n16, A2 => net31039, A3 => n15, ZN => p(3));
   U52 : MUX2_X1 port map( A => net31025, B => net31021, S => A(3), Z => n18);
   U53 : MUX2_X1 port map( A => n7, B => net31045, S => A(4), Z => n17);
   U54 : NAND3_X1 port map( A1 => n18, A2 => net31039, A3 => n17, ZN => p(4));
   U55 : MUX2_X1 port map( A => n7, B => n2, S => A(5), Z => n20);
   U56 : MUX2_X1 port map( A => net31027, B => net31021, S => A(4), Z => n19);
   U57 : NAND3_X1 port map( A1 => n20, A2 => net31039, A3 => n19, ZN => p(5));
   U58 : MUX2_X1 port map( A => net31029, B => net31021, S => A(5), Z => n22);
   U59 : MUX2_X1 port map( A => net31033, B => net31045, S => A(6), Z => n21);
   U60 : NAND3_X1 port map( A1 => n22, A2 => net31039, A3 => n21, ZN => p(6));
   U61 : MUX2_X1 port map( A => net31027, B => net31021, S => A(6), Z => n24);
   U62 : MUX2_X1 port map( A => net31031, B => n2, S => A(7), Z => n23);
   U63 : NAND3_X1 port map( A1 => n24, A2 => net31039, A3 => n23, ZN => p(7));
   U64 : MUX2_X1 port map( A => net31029, B => net31021, S => A(7), Z => n26);
   U65 : MUX2_X1 port map( A => net31031, B => net31045, S => A(8), Z => n25);
   U66 : NAND3_X1 port map( A1 => n26, A2 => net31037, A3 => n25, ZN => p(8));
   U67 : MUX2_X1 port map( A => net31027, B => net31021, S => A(8), Z => n28);
   U68 : MUX2_X1 port map( A => n7, B => net31045, S => A(9), Z => n27);
   U69 : NAND3_X1 port map( A1 => n28, A2 => net31037, A3 => n27, ZN => p(9));
   U70 : MUX2_X1 port map( A => net31027, B => net31021, S => A(9), Z => n32);
   U71 : XOR2_X1 port map( A => b(1), B => b(0), Z => n29);
   U72 : NAND2_X1 port map( A1 => n29, A2 => net29502, ZN => n30);
   U73 : MUX2_X1 port map( A => n7, B => n30, S => A(10), Z => n31);
   U74 : NAND3_X1 port map( A1 => n32, A2 => net31037, A3 => n31, ZN => p(10));
   U75 : MUX2_X1 port map( A => net31029, B => net31021, S => A(10), Z => n34);
   U76 : MUX2_X1 port map( A => n7, B => net31045, S => A(11), Z => n33);
   U77 : NAND3_X1 port map( A1 => n34, A2 => net31037, A3 => n33, ZN => p(11));
   U78 : MUX2_X1 port map( A => net31027, B => net31021, S => A(11), Z => n36);
   U79 : MUX2_X1 port map( A => net31033, B => net31045, S => A(12), Z => n35);
   U80 : NAND3_X1 port map( A1 => n36, A2 => net31037, A3 => n35, ZN => p(12));
   U81 : MUX2_X1 port map( A => net31025, B => net31021, S => A(12), Z => n37);
   U82 : NAND3_X1 port map( A1 => net29492, A2 => n37, A3 => net31037, ZN => 
                           p(13));
   U83 : MUX2_X1 port map( A => net31031, B => net31045, S => A(15), Z => n38);
   U84 : NAND3_X1 port map( A1 => net29488, A2 => net31037, A3 => n38, ZN => 
                           p(15));
   U85 : MUX2_X1 port map( A => net31027, B => net31021, S => A(15), Z => n40);
   U86 : MUX2_X1 port map( A => net31033, B => net31045, S => A(16), Z => n39);
   U87 : NAND3_X1 port map( A1 => n40, A2 => net31037, A3 => n39, ZN => p(16));
   U88 : MUX2_X1 port map( A => net31029, B => net31021, S => A(16), Z => n42);
   U89 : MUX2_X1 port map( A => net31033, B => net31045, S => A(17), Z => n41);
   U90 : NAND3_X1 port map( A1 => n42, A2 => net31037, A3 => n41, ZN => p(17));
   U91 : MUX2_X1 port map( A => net31029, B => net31019, S => A(17), Z => n44);
   U92 : MUX2_X1 port map( A => net31031, B => net31045, S => A(18), Z => n43);
   U93 : NAND3_X1 port map( A1 => n44, A2 => net31037, A3 => n43, ZN => p(18));
   U94 : MUX2_X1 port map( A => n7, B => n2, S => A(19), Z => n46);
   U95 : MUX2_X1 port map( A => net31025, B => net31019, S => A(18), Z => n45);
   U96 : NAND3_X1 port map( A1 => net31039, A2 => n46, A3 => n45, ZN => p(19));
   U97 : MUX2_X1 port map( A => net31029, B => net31019, S => A(19), Z => n48);
   U98 : MUX2_X1 port map( A => net31031, B => n2, S => A(20), Z => n47);
   U99 : NAND3_X1 port map( A1 => n48, A2 => net31035, A3 => n47, ZN => p(20));
   U100 : MUX2_X1 port map( A => net31027, B => net31019, S => A(20), Z => n50)
                           ;
   U101 : MUX2_X1 port map( A => net31031, B => net31045, S => A(21), Z => n49)
                           ;
   U102 : NAND3_X1 port map( A1 => n50, A2 => net31037, A3 => n49, ZN => p(21))
                           ;
   U103 : MUX2_X1 port map( A => net31027, B => net31019, S => A(21), Z => n52)
                           ;
   U104 : MUX2_X1 port map( A => n7, B => n2, S => A(22), Z => n51);
   U105 : NAND3_X1 port map( A1 => n52, A2 => net31035, A3 => n51, ZN => p(22))
                           ;
   U106 : MUX2_X1 port map( A => net31029, B => net31019, S => A(22), Z => n54)
                           ;
   U107 : MUX2_X1 port map( A => n7, B => n2, S => A(23), Z => n53);
   U108 : NAND3_X1 port map( A1 => n54, A2 => net31035, A3 => n53, ZN => p(23))
                           ;
   U109 : MUX2_X1 port map( A => net31029, B => net31019, S => A(23), Z => n56)
                           ;
   U110 : MUX2_X1 port map( A => net31033, B => n2, S => A(24), Z => n55);
   U111 : NAND3_X1 port map( A1 => n56, A2 => net31035, A3 => n55, ZN => p(24))
                           ;
   U112 : MUX2_X1 port map( A => net31029, B => net31019, S => A(24), Z => n58)
                           ;
   U113 : MUX2_X1 port map( A => net31033, B => n2, S => A(25), Z => n57);
   U114 : NAND3_X1 port map( A1 => n58, A2 => net31035, A3 => n57, ZN => p(25))
                           ;
   U115 : MUX2_X1 port map( A => net31031, B => net31045, S => A(26), Z => n59)
                           ;
   U116 : NAND3_X1 port map( A1 => n60, A2 => net31035, A3 => n59, ZN => p(26))
                           ;
   U117 : MUX2_X1 port map( A => net31033, B => n2, S => A(27), Z => n61);
   U118 : NAND3_X1 port map( A1 => n62, A2 => net31035, A3 => n61, ZN => p(27))
                           ;
   U119 : MUX2_X1 port map( A => n7, B => n2, S => A(28), Z => n63);
   U120 : NAND3_X1 port map( A1 => n64, A2 => net31035, A3 => n63, ZN => p(28))
                           ;
   U121 : MUX2_X1 port map( A => net31031, B => net31045, S => A(29), Z => n65)
                           ;
   U122 : NAND3_X1 port map( A1 => n66, A2 => net31035, A3 => n65, ZN => p(29))
                           ;
   U123 : MUX2_X1 port map( A => net31033, B => n1, S => A(30), Z => n67);
   U124 : NAND3_X1 port map( A1 => n68, A2 => net31035, A3 => n67, ZN => p(30))
                           ;
   U125 : MUX2_X1 port map( A => n7, B => n1, S => n8, Z => n69);
   U126 : NAND3_X1 port map( A1 => n70, A2 => net31035, A3 => n69, ZN => p(31))
                           ;
   U127 : OAI221_X1 port map( B1 => n9, B2 => net31019, C1 => n8, C2 => 
                           net31027, A => net31031, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_5 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_5;

architecture SYN_beh of ENC_5 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90 : std_logic;

begin
   
   U3 : OR2_X1 port map( A1 => b(2), A2 => n16, ZN => n84);
   U4 : CLKBUF_X3 port map( A => n86, Z => n5);
   U5 : CLKBUF_X3 port map( A => n86, Z => n4);
   U6 : BUF_X1 port map( A => n84, Z => n2);
   U7 : BUF_X2 port map( A => n84, Z => n1);
   U8 : BUF_X1 port map( A => n88, Z => n7);
   U9 : BUF_X1 port map( A => n90, Z => n13);
   U10 : BUF_X1 port map( A => n89, Z => n10);
   U11 : BUF_X1 port map( A => n88, Z => n8);
   U12 : MUX2_X1 port map( A => n10, B => n12, S => A(28), Z => n81);
   U13 : MUX2_X1 port map( A => n11, B => n12, S => A(29), Z => n83);
   U14 : MUX2_X1 port map( A => n10, B => n12, S => A(27), Z => n79);
   U15 : BUF_X1 port map( A => n90, Z => n12);
   U16 : BUF_X1 port map( A => n89, Z => n9);
   U17 : MUX2_X1 port map( A => n10, B => n12, S => A(24), Z => n73);
   U18 : MUX2_X1 port map( A => n10, B => n12, S => A(25), Z => n75);
   U19 : MUX2_X1 port map( A => n10, B => n12, S => A(26), Z => n77);
   U20 : MUX2_X1 port map( A => n10, B => n12, S => A(23), Z => n71);
   U21 : MUX2_X1 port map( A => n11, B => n12, S => A(30), Z => n87);
   U22 : CLKBUF_X1 port map( A => n84, Z => n3);
   U23 : BUF_X1 port map( A => n90, Z => n14);
   U24 : BUF_X1 port map( A => n89, Z => n11);
   U25 : XNOR2_X1 port map( A => b(1), B => b(0), ZN => n16);
   U26 : BUF_X2 port map( A => n86, Z => n6);
   U27 : INV_X1 port map( A => A(31), ZN => n15);
   U28 : INV_X1 port map( A => b(2), ZN => n19);
   U29 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n18);
   U30 : INV_X1 port map( A => b(0), ZN => n21);
   U31 : INV_X1 port map( A => b(1), ZN => n20);
   U32 : NAND3_X1 port map( A1 => b(2), A2 => n21, A3 => n20, ZN => n89);
   U33 : NAND2_X1 port map( A1 => b(2), A2 => n18, ZN => n22);
   U34 : MUX2_X1 port map( A => n22, B => n2, S => A(0), Z => n17);
   U35 : OAI211_X1 port map( C1 => n19, C2 => n18, A => n9, B => n17, ZN => 
                           p(0));
   U36 : NAND3_X1 port map( A1 => b(1), A2 => n19, A3 => b(0), ZN => n90);
   U37 : MUX2_X1 port map( A => n9, B => n13, S => A(0), Z => n25);
   U38 : NAND2_X1 port map( A1 => n21, A2 => n20, ZN => n23);
   U39 : NAND4_X1 port map( A1 => n1, A2 => n22, A3 => n23, A4 => n12, ZN => 
                           n86);
   U40 : NAND2_X1 port map( A1 => b(2), A2 => n23, ZN => n88);
   U41 : MUX2_X1 port map( A => n8, B => n1, S => A(1), Z => n24);
   U42 : NAND3_X1 port map( A1 => n25, A2 => n4, A3 => n24, ZN => p(1));
   U43 : MUX2_X1 port map( A => n8, B => n1, S => A(2), Z => n27);
   U44 : MUX2_X1 port map( A => n9, B => n12, S => A(1), Z => n26);
   U45 : NAND3_X1 port map( A1 => n27, A2 => n26, A3 => n4, ZN => p(2));
   U46 : MUX2_X1 port map( A => n9, B => n12, S => A(2), Z => n29);
   U47 : MUX2_X1 port map( A => n8, B => n1, S => A(3), Z => n28);
   U48 : NAND3_X1 port map( A1 => n29, A2 => n6, A3 => n28, ZN => p(3));
   U49 : MUX2_X1 port map( A => n9, B => n12, S => A(3), Z => n31);
   U50 : MUX2_X1 port map( A => n8, B => n1, S => A(4), Z => n30);
   U51 : NAND3_X1 port map( A1 => n31, A2 => n6, A3 => n30, ZN => p(4));
   U52 : MUX2_X1 port map( A => n8, B => n1, S => A(5), Z => n33);
   U53 : MUX2_X1 port map( A => n9, B => n12, S => A(4), Z => n32);
   U54 : NAND3_X1 port map( A1 => n33, A2 => n6, A3 => n32, ZN => p(5));
   U55 : MUX2_X1 port map( A => n8, B => n1, S => A(6), Z => n35);
   U56 : MUX2_X1 port map( A => n9, B => n13, S => A(5), Z => n34);
   U57 : NAND3_X1 port map( A1 => n35, A2 => n6, A3 => n34, ZN => p(6));
   U58 : MUX2_X1 port map( A => n8, B => n1, S => A(7), Z => n37);
   U59 : MUX2_X1 port map( A => n9, B => n13, S => A(6), Z => n36);
   U60 : NAND3_X1 port map( A1 => n6, A2 => n37, A3 => n36, ZN => p(7));
   U61 : MUX2_X1 port map( A => n9, B => n13, S => A(7), Z => n39);
   U62 : MUX2_X1 port map( A => n8, B => n1, S => A(8), Z => n38);
   U63 : NAND3_X1 port map( A1 => n39, A2 => n6, A3 => n38, ZN => p(8));
   U64 : MUX2_X1 port map( A => n10, B => n13, S => A(8), Z => n41);
   U65 : MUX2_X1 port map( A => n8, B => n1, S => A(9), Z => n40);
   U66 : NAND3_X1 port map( A1 => n41, A2 => n6, A3 => n40, ZN => p(9));
   U67 : MUX2_X1 port map( A => n9, B => n13, S => A(9), Z => n43);
   U68 : MUX2_X1 port map( A => n8, B => n1, S => A(10), Z => n42);
   U69 : NAND3_X1 port map( A1 => n43, A2 => n5, A3 => n42, ZN => p(10));
   U70 : MUX2_X1 port map( A => n9, B => n13, S => A(10), Z => n45);
   U71 : MUX2_X1 port map( A => n8, B => n1, S => A(11), Z => n44);
   U72 : NAND3_X1 port map( A1 => n45, A2 => n5, A3 => n44, ZN => p(11));
   U73 : MUX2_X1 port map( A => n9, B => n13, S => A(11), Z => n47);
   U74 : MUX2_X1 port map( A => n8, B => n1, S => A(12), Z => n46);
   U75 : NAND3_X1 port map( A1 => n47, A2 => n5, A3 => n46, ZN => p(12));
   U76 : MUX2_X1 port map( A => n9, B => n13, S => A(12), Z => n49);
   U77 : MUX2_X1 port map( A => n8, B => n1, S => A(13), Z => n48);
   U78 : NAND3_X1 port map( A1 => n49, A2 => n5, A3 => n48, ZN => p(13));
   U79 : MUX2_X1 port map( A => n9, B => n13, S => A(13), Z => n51);
   U80 : MUX2_X1 port map( A => n8, B => n2, S => A(14), Z => n50);
   U81 : NAND3_X1 port map( A1 => n51, A2 => n5, A3 => n50, ZN => p(14));
   U82 : MUX2_X1 port map( A => n10, B => n13, S => A(14), Z => n53);
   U83 : MUX2_X1 port map( A => n8, B => n2, S => A(15), Z => n52);
   U84 : NAND3_X1 port map( A1 => n53, A2 => n5, A3 => n52, ZN => p(15));
   U85 : MUX2_X1 port map( A => n10, B => n13, S => A(15), Z => n55);
   U86 : MUX2_X1 port map( A => n8, B => n2, S => A(16), Z => n54);
   U87 : NAND3_X1 port map( A1 => n55, A2 => n5, A3 => n54, ZN => p(16));
   U88 : MUX2_X1 port map( A => n10, B => n13, S => A(16), Z => n57);
   U89 : MUX2_X1 port map( A => n7, B => n2, S => A(17), Z => n56);
   U90 : NAND3_X1 port map( A1 => n57, A2 => n5, A3 => n56, ZN => p(17));
   U91 : MUX2_X1 port map( A => n10, B => n13, S => A(17), Z => n59);
   U92 : MUX2_X1 port map( A => n7, B => n2, S => A(18), Z => n58);
   U93 : NAND3_X1 port map( A1 => n59, A2 => n5, A3 => n58, ZN => p(18));
   U94 : MUX2_X1 port map( A => n10, B => n13, S => A(18), Z => n61);
   U95 : MUX2_X1 port map( A => n7, B => n2, S => A(19), Z => n60);
   U96 : NAND3_X1 port map( A1 => n61, A2 => n5, A3 => n60, ZN => p(19));
   U97 : MUX2_X1 port map( A => n10, B => n13, S => A(19), Z => n63);
   U98 : MUX2_X1 port map( A => n7, B => n2, S => A(20), Z => n62);
   U99 : NAND3_X1 port map( A1 => n63, A2 => n5, A3 => n62, ZN => p(20));
   U100 : MUX2_X1 port map( A => n10, B => n14, S => A(20), Z => n65);
   U101 : MUX2_X1 port map( A => n7, B => n2, S => A(21), Z => n64);
   U102 : NAND3_X1 port map( A1 => n65, A2 => n4, A3 => n64, ZN => p(21));
   U103 : MUX2_X1 port map( A => n10, B => n14, S => A(21), Z => n67);
   U104 : MUX2_X1 port map( A => n7, B => n2, S => A(22), Z => n66);
   U105 : NAND3_X1 port map( A1 => n67, A2 => n4, A3 => n66, ZN => p(22));
   U106 : MUX2_X1 port map( A => n10, B => n12, S => A(22), Z => n69);
   U107 : MUX2_X1 port map( A => n7, B => n2, S => A(23), Z => n68);
   U108 : NAND3_X1 port map( A1 => n69, A2 => n4, A3 => n68, ZN => p(23));
   U109 : MUX2_X1 port map( A => n7, B => n2, S => A(24), Z => n70);
   U110 : NAND3_X1 port map( A1 => n71, A2 => n4, A3 => n70, ZN => p(24));
   U111 : MUX2_X1 port map( A => n7, B => n2, S => A(25), Z => n72);
   U112 : NAND3_X1 port map( A1 => n73, A2 => n4, A3 => n72, ZN => p(25));
   U113 : MUX2_X1 port map( A => n7, B => n2, S => A(26), Z => n74);
   U114 : NAND3_X1 port map( A1 => n75, A2 => n4, A3 => n74, ZN => p(26));
   U115 : MUX2_X1 port map( A => n7, B => n2, S => A(27), Z => n76);
   U116 : NAND3_X1 port map( A1 => n77, A2 => n4, A3 => n76, ZN => p(27));
   U117 : MUX2_X1 port map( A => n7, B => n3, S => A(28), Z => n78);
   U118 : NAND3_X1 port map( A1 => n79, A2 => n4, A3 => n78, ZN => p(28));
   U119 : MUX2_X1 port map( A => n7, B => n3, S => A(29), Z => n80);
   U120 : NAND3_X1 port map( A1 => n81, A2 => n4, A3 => n80, ZN => p(29));
   U121 : MUX2_X1 port map( A => n7, B => n3, S => A(30), Z => n82);
   U122 : NAND3_X1 port map( A1 => n83, A2 => n4, A3 => n82, ZN => p(30));
   U123 : MUX2_X1 port map( A => n7, B => n1, S => A(31), Z => n85);
   U124 : NAND3_X1 port map( A1 => n87, A2 => n5, A3 => n85, ZN => p(31));
   U125 : OAI221_X1 port map( B1 => n15, B2 => n12, C1 => A(31), C2 => n9, A =>
                           n7, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_4 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_4;

architecture SYN_beh of ENC_4 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95 : std_logic;

begin
   
   U3 : BUF_X1 port map( A => n91, Z => n4);
   U4 : BUF_X1 port map( A => n91, Z => n5);
   U5 : INV_X1 port map( A => n7, ZN => n6);
   U6 : MUX2_X1 port map( A => n9, B => n11, S => A(22), Z => n74);
   U7 : MUX2_X1 port map( A => n9, B => n11, S => A(23), Z => n76);
   U8 : MUX2_X1 port map( A => n9, B => n11, S => A(21), Z => n72);
   U9 : BUF_X1 port map( A => n95, Z => n11);
   U10 : BUF_X1 port map( A => n94, Z => n9);
   U11 : BUF_X1 port map( A => n95, Z => n12);
   U12 : BUF_X1 port map( A => n94, Z => n8);
   U13 : BUF_X1 port map( A => n89, Z => n1);
   U14 : BUF_X1 port map( A => n89, Z => n2);
   U15 : BUF_X1 port map( A => n89, Z => n3);
   U16 : BUF_X1 port map( A => n95, Z => n13);
   U17 : BUF_X1 port map( A => n94, Z => n10);
   U18 : INV_X1 port map( A => n93, ZN => n7);
   U19 : INV_X1 port map( A => A(24), ZN => n14);
   U20 : INV_X1 port map( A => A(25), ZN => n15);
   U21 : INV_X1 port map( A => A(26), ZN => n16);
   U22 : INV_X1 port map( A => A(27), ZN => n17);
   U23 : INV_X1 port map( A => A(28), ZN => n18);
   U24 : INV_X1 port map( A => A(29), ZN => n19);
   U25 : INV_X1 port map( A => A(30), ZN => n20);
   U26 : INV_X1 port map( A => A(31), ZN => n21);
   U27 : INV_X1 port map( A => b(2), ZN => n26);
   U28 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n95);
   U29 : INV_X1 port map( A => b(0), ZN => n23);
   U30 : INV_X1 port map( A => b(1), ZN => n22);
   U31 : NAND3_X1 port map( A1 => b(2), A2 => n23, A3 => n22, ZN => n94);
   U32 : NAND2_X1 port map( A1 => b(2), A2 => n11, ZN => n31);
   U33 : XOR2_X1 port map( A => b(1), B => b(0), Z => n24);
   U34 : NAND2_X1 port map( A1 => n24, A2 => n26, ZN => n89);
   U35 : MUX2_X1 port map( A => n31, B => n3, S => A(0), Z => n25);
   U36 : OAI211_X1 port map( C1 => n26, C2 => n11, A => n8, B => n25, ZN => 
                           p(0));
   U37 : MUX2_X1 port map( A => n8, B => n11, S => A(0), Z => n28);
   U38 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => b(2), ZN => n93);
   U39 : NAND2_X1 port map( A1 => n7, A2 => n31, ZN => n91);
   U40 : MUX2_X1 port map( A => n93, B => n3, S => A(1), Z => n27);
   U41 : NAND3_X1 port map( A1 => n28, A2 => n5, A3 => n27, ZN => p(1));
   U42 : MUX2_X1 port map( A => n93, B => n3, S => A(2), Z => n30);
   U43 : MUX2_X1 port map( A => n8, B => n12, S => A(1), Z => n29);
   U44 : NAND3_X1 port map( A1 => n30, A2 => n29, A3 => n4, ZN => p(2));
   U45 : MUX2_X1 port map( A => n8, B => n12, S => A(2), Z => n33);
   U46 : NAND2_X1 port map( A1 => n7, A2 => n31, ZN => n51);
   U47 : MUX2_X1 port map( A => n93, B => n3, S => A(3), Z => n32);
   U48 : NAND3_X1 port map( A1 => n33, A2 => n51, A3 => n32, ZN => p(3));
   U49 : MUX2_X1 port map( A => n8, B => n12, S => A(3), Z => n35);
   U50 : MUX2_X1 port map( A => n93, B => n3, S => A(4), Z => n34);
   U51 : NAND3_X1 port map( A1 => n35, A2 => n51, A3 => n34, ZN => p(4));
   U52 : MUX2_X1 port map( A => n93, B => n3, S => A(5), Z => n37);
   U53 : MUX2_X1 port map( A => n8, B => n12, S => A(4), Z => n36);
   U54 : NAND3_X1 port map( A1 => n37, A2 => n36, A3 => n51, ZN => p(5));
   U55 : MUX2_X1 port map( A => n8, B => n12, S => A(5), Z => n39);
   U56 : MUX2_X1 port map( A => n93, B => n3, S => A(6), Z => n38);
   U57 : NAND3_X1 port map( A1 => n39, A2 => n51, A3 => n38, ZN => p(6));
   U58 : MUX2_X1 port map( A => n8, B => n12, S => A(6), Z => n41);
   U59 : MUX2_X1 port map( A => n93, B => n3, S => A(7), Z => n40);
   U60 : NAND3_X1 port map( A1 => n41, A2 => n51, A3 => n40, ZN => p(7));
   U61 : MUX2_X1 port map( A => n8, B => n12, S => A(7), Z => n43);
   U62 : MUX2_X1 port map( A => n93, B => n3, S => A(8), Z => n42);
   U63 : NAND3_X1 port map( A1 => n43, A2 => n4, A3 => n42, ZN => p(8));
   U64 : MUX2_X1 port map( A => n9, B => n12, S => A(8), Z => n45);
   U65 : MUX2_X1 port map( A => n93, B => n3, S => A(9), Z => n44);
   U66 : NAND3_X1 port map( A1 => n45, A2 => n4, A3 => n44, ZN => p(9));
   U67 : MUX2_X1 port map( A => n8, B => n12, S => A(9), Z => n47);
   U68 : MUX2_X1 port map( A => n93, B => n2, S => A(10), Z => n46);
   U69 : NAND3_X1 port map( A1 => n47, A2 => n4, A3 => n46, ZN => p(10));
   U70 : MUX2_X1 port map( A => n8, B => n12, S => A(10), Z => n49);
   U71 : MUX2_X1 port map( A => n93, B => n2, S => A(11), Z => n48);
   U72 : NAND3_X1 port map( A1 => n49, A2 => n4, A3 => n48, ZN => p(11));
   U73 : MUX2_X1 port map( A => n8, B => n12, S => A(11), Z => n52);
   U74 : MUX2_X1 port map( A => n93, B => n2, S => A(12), Z => n50);
   U75 : NAND3_X1 port map( A1 => n52, A2 => n51, A3 => n50, ZN => p(12));
   U76 : MUX2_X1 port map( A => n8, B => n12, S => A(12), Z => n54);
   U77 : MUX2_X1 port map( A => n93, B => n2, S => A(13), Z => n53);
   U78 : NAND3_X1 port map( A1 => n54, A2 => n4, A3 => n53, ZN => p(13));
   U79 : MUX2_X1 port map( A => n8, B => n12, S => A(13), Z => n56);
   U80 : MUX2_X1 port map( A => n93, B => n2, S => A(14), Z => n55);
   U81 : NAND3_X1 port map( A1 => n56, A2 => n4, A3 => n55, ZN => p(14));
   U82 : MUX2_X1 port map( A => n9, B => n12, S => A(14), Z => n58);
   U83 : MUX2_X1 port map( A => n93, B => n2, S => A(15), Z => n57);
   U84 : NAND3_X1 port map( A1 => n58, A2 => n4, A3 => n57, ZN => p(15));
   U85 : MUX2_X1 port map( A => n6, B => n2, S => A(16), Z => n60);
   U86 : MUX2_X1 port map( A => n9, B => n12, S => A(15), Z => n59);
   U87 : NAND3_X1 port map( A1 => n91, A2 => n60, A3 => n59, ZN => p(16));
   U88 : MUX2_X1 port map( A => n9, B => n12, S => A(16), Z => n62);
   U89 : MUX2_X1 port map( A => n6, B => n2, S => A(17), Z => n61);
   U90 : NAND3_X1 port map( A1 => n62, A2 => n4, A3 => n61, ZN => p(17));
   U91 : MUX2_X1 port map( A => n9, B => n13, S => A(17), Z => n64);
   U92 : MUX2_X1 port map( A => n6, B => n2, S => A(18), Z => n63);
   U93 : NAND3_X1 port map( A1 => n64, A2 => n4, A3 => n63, ZN => p(18));
   U94 : MUX2_X1 port map( A => n9, B => n13, S => A(18), Z => n66);
   U95 : MUX2_X1 port map( A => n6, B => n2, S => A(19), Z => n65);
   U96 : NAND3_X1 port map( A1 => n66, A2 => n4, A3 => n65, ZN => p(19));
   U97 : MUX2_X1 port map( A => n9, B => n13, S => A(19), Z => n68);
   U98 : MUX2_X1 port map( A => n6, B => n2, S => A(20), Z => n67);
   U99 : NAND3_X1 port map( A1 => n68, A2 => n5, A3 => n67, ZN => p(20));
   U100 : MUX2_X1 port map( A => n9, B => n11, S => A(20), Z => n70);
   U101 : MUX2_X1 port map( A => n6, B => n1, S => A(21), Z => n69);
   U102 : NAND3_X1 port map( A1 => n70, A2 => n5, A3 => n69, ZN => p(21));
   U103 : MUX2_X1 port map( A => n6, B => n1, S => A(22), Z => n71);
   U104 : NAND3_X1 port map( A1 => n72, A2 => n5, A3 => n71, ZN => p(22));
   U105 : MUX2_X1 port map( A => n6, B => n1, S => A(23), Z => n73);
   U106 : NAND3_X1 port map( A1 => n74, A2 => n5, A3 => n73, ZN => p(23));
   U107 : MUX2_X1 port map( A => n6, B => n1, S => A(24), Z => n75);
   U108 : NAND3_X1 port map( A1 => n76, A2 => n5, A3 => n75, ZN => p(24));
   U109 : MUX2_X1 port map( A => n11, B => n9, S => n14, Z => n78);
   U110 : MUX2_X1 port map( A => n6, B => n1, S => A(25), Z => n77);
   U111 : NAND3_X1 port map( A1 => n78, A2 => n5, A3 => n77, ZN => p(25));
   U112 : MUX2_X1 port map( A => n11, B => n9, S => n15, Z => n80);
   U113 : MUX2_X1 port map( A => n6, B => n1, S => A(26), Z => n79);
   U114 : NAND3_X1 port map( A1 => n80, A2 => n5, A3 => n79, ZN => p(26));
   U115 : MUX2_X1 port map( A => n11, B => n9, S => n16, Z => n82);
   U116 : MUX2_X1 port map( A => n6, B => n1, S => A(27), Z => n81);
   U117 : NAND3_X1 port map( A1 => n82, A2 => n5, A3 => n81, ZN => p(27));
   U118 : MUX2_X1 port map( A => n11, B => n9, S => n17, Z => n84);
   U119 : MUX2_X1 port map( A => n6, B => n1, S => A(28), Z => n83);
   U120 : NAND3_X1 port map( A1 => n84, A2 => n5, A3 => n83, ZN => p(28));
   U121 : MUX2_X1 port map( A => n11, B => n9, S => n18, Z => n86);
   U122 : MUX2_X1 port map( A => n6, B => n1, S => A(29), Z => n85);
   U123 : NAND3_X1 port map( A1 => n86, A2 => n5, A3 => n85, ZN => p(29));
   U124 : MUX2_X1 port map( A => n11, B => n10, S => n19, Z => n88);
   U125 : MUX2_X1 port map( A => n6, B => n1, S => A(30), Z => n87);
   U126 : NAND3_X1 port map( A1 => n88, A2 => n5, A3 => n87, ZN => p(30));
   U127 : MUX2_X1 port map( A => n11, B => n10, S => n20, Z => n92);
   U128 : MUX2_X1 port map( A => n6, B => n1, S => A(31), Z => n90);
   U129 : NAND3_X1 port map( A1 => n92, A2 => n4, A3 => n90, ZN => p(31));
   U130 : OAI221_X1 port map( B1 => n21, B2 => n11, C1 => A(31), C2 => n8, A =>
                           n6, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_3 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_3;

architecture SYN_beh of ENC_3 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   U3 : BUF_X1 port map( A => n95, Z => n6);
   U4 : BUF_X1 port map( A => n95, Z => n7);
   U5 : BUF_X1 port map( A => n95, Z => n8);
   U6 : BUF_X1 port map( A => n97, Z => n9);
   U7 : MUX2_X1 port map( A => n12, B => n14, S => A(21), Z => n76);
   U8 : MUX2_X1 port map( A => n12, B => n14, S => A(20), Z => n74);
   U9 : MUX2_X1 port map( A => n12, B => n14, S => A(22), Z => n78);
   U10 : MUX2_X1 port map( A => n12, B => n14, S => A(19), Z => n72);
   U11 : MUX2_X1 port map( A => n12, B => n14, S => A(23), Z => n80);
   U12 : BUF_X1 port map( A => n98, Z => n12);
   U13 : BUF_X1 port map( A => n98, Z => n11);
   U14 : BUF_X1 port map( A => n99, Z => n14);
   U15 : BUF_X1 port map( A => n97, Z => n10);
   U16 : BUF_X1 port map( A => n99, Z => n15);
   U17 : BUF_X1 port map( A => n93, Z => n3);
   U18 : BUF_X1 port map( A => n93, Z => n4);
   U19 : BUF_X1 port map( A => n93, Z => n5);
   U20 : BUF_X1 port map( A => n98, Z => n13);
   U21 : OR2_X1 port map( A1 => b(2), A2 => n22, ZN => n93);
   U22 : XNOR2_X1 port map( A => b(1), B => b(0), ZN => n22);
   U23 : INV_X1 port map( A => A(29), ZN => n1);
   U24 : INV_X1 port map( A => A(30), ZN => n2);
   U25 : INV_X1 port map( A => A(24), ZN => n16);
   U26 : INV_X1 port map( A => A(25), ZN => n17);
   U27 : INV_X1 port map( A => A(26), ZN => n18);
   U28 : INV_X1 port map( A => A(27), ZN => n19);
   U29 : INV_X1 port map( A => A(28), ZN => n20);
   U30 : INV_X1 port map( A => A(31), ZN => n21);
   U31 : INV_X1 port map( A => b(2), ZN => n25);
   U32 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n24);
   U33 : INV_X1 port map( A => b(0), ZN => n27);
   U34 : INV_X1 port map( A => b(1), ZN => n26);
   U35 : NAND3_X1 port map( A1 => b(2), A2 => n27, A3 => n26, ZN => n98);
   U36 : NAND2_X1 port map( A1 => b(2), A2 => n24, ZN => n28);
   U37 : MUX2_X1 port map( A => n28, B => n5, S => A(0), Z => n23);
   U38 : OAI211_X1 port map( C1 => n25, C2 => n24, A => n11, B => n23, ZN => 
                           p(0));
   U39 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n99);
   U40 : MUX2_X1 port map( A => n11, B => n15, S => A(0), Z => n32);
   U41 : NAND2_X1 port map( A1 => n27, A2 => n26, ZN => n30);
   U42 : NAND2_X1 port map( A1 => b(2), A2 => n30, ZN => n39);
   U43 : INV_X1 port map( A => n39, ZN => n29);
   U44 : NAND2_X1 port map( A1 => n29, A2 => n28, ZN => n95);
   U45 : NAND2_X1 port map( A1 => b(2), A2 => n30, ZN => n97);
   U46 : MUX2_X1 port map( A => n10, B => n5, S => A(1), Z => n31);
   U47 : NAND3_X1 port map( A1 => n32, A2 => n6, A3 => n31, ZN => p(1));
   U48 : MUX2_X1 port map( A => n11, B => n15, S => A(1), Z => n34);
   U49 : MUX2_X1 port map( A => n39, B => n5, S => A(2), Z => n33);
   U50 : NAND3_X1 port map( A1 => n34, A2 => n8, A3 => n33, ZN => p(2));
   U51 : MUX2_X1 port map( A => n11, B => n15, S => A(2), Z => n36);
   U52 : MUX2_X1 port map( A => n39, B => n5, S => A(3), Z => n35);
   U53 : NAND3_X1 port map( A1 => n36, A2 => n8, A3 => n35, ZN => p(3));
   U54 : MUX2_X1 port map( A => n39, B => n5, S => A(4), Z => n38);
   U55 : MUX2_X1 port map( A => n11, B => n15, S => A(3), Z => n37);
   U56 : NAND3_X1 port map( A1 => n38, A2 => n37, A3 => n6, ZN => p(4));
   U57 : MUX2_X1 port map( A => n39, B => n5, S => A(5), Z => n41);
   U58 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n60);
   U59 : MUX2_X1 port map( A => n11, B => n60, S => A(4), Z => n40);
   U60 : NAND3_X1 port map( A1 => n41, A2 => n40, A3 => n6, ZN => p(5));
   U61 : MUX2_X1 port map( A => n11, B => n15, S => A(5), Z => n43);
   U62 : MUX2_X1 port map( A => n10, B => n5, S => A(6), Z => n42);
   U63 : NAND3_X1 port map( A1 => n43, A2 => n8, A3 => n42, ZN => p(6));
   U64 : MUX2_X1 port map( A => n11, B => n15, S => A(6), Z => n45);
   U65 : MUX2_X1 port map( A => n10, B => n5, S => A(7), Z => n44);
   U66 : NAND3_X1 port map( A1 => n45, A2 => n8, A3 => n44, ZN => p(7));
   U67 : MUX2_X1 port map( A => n11, B => n15, S => A(7), Z => n47);
   U68 : MUX2_X1 port map( A => n10, B => n5, S => A(8), Z => n46);
   U69 : NAND3_X1 port map( A1 => n47, A2 => n8, A3 => n46, ZN => p(8));
   U70 : MUX2_X1 port map( A => n12, B => n15, S => A(8), Z => n49);
   U71 : MUX2_X1 port map( A => n10, B => n5, S => A(9), Z => n48);
   U72 : NAND3_X1 port map( A1 => n49, A2 => n8, A3 => n48, ZN => p(9));
   U73 : MUX2_X1 port map( A => n11, B => n60, S => A(9), Z => n51);
   U74 : MUX2_X1 port map( A => n10, B => n4, S => A(10), Z => n50);
   U75 : NAND3_X1 port map( A1 => n51, A2 => n7, A3 => n50, ZN => p(10));
   U76 : MUX2_X1 port map( A => n11, B => n60, S => A(10), Z => n53);
   U77 : MUX2_X1 port map( A => n10, B => n4, S => A(11), Z => n52);
   U78 : NAND3_X1 port map( A1 => n53, A2 => n7, A3 => n52, ZN => p(11));
   U79 : MUX2_X1 port map( A => n10, B => n4, S => A(12), Z => n55);
   U80 : MUX2_X1 port map( A => n11, B => n60, S => A(11), Z => n54);
   U81 : NAND3_X1 port map( A1 => n55, A2 => n54, A3 => n6, ZN => p(12));
   U82 : MUX2_X1 port map( A => n11, B => n15, S => A(12), Z => n57);
   U83 : MUX2_X1 port map( A => n10, B => n4, S => A(13), Z => n56);
   U84 : NAND3_X1 port map( A1 => n57, A2 => n7, A3 => n56, ZN => p(13));
   U85 : MUX2_X1 port map( A => n10, B => n4, S => A(14), Z => n59);
   U86 : MUX2_X1 port map( A => n11, B => n15, S => A(13), Z => n58);
   U87 : NAND3_X1 port map( A1 => n8, A2 => n59, A3 => n58, ZN => p(14));
   U88 : MUX2_X1 port map( A => n12, B => n60, S => A(14), Z => n62);
   U89 : MUX2_X1 port map( A => n10, B => n4, S => A(15), Z => n61);
   U90 : NAND3_X1 port map( A1 => n62, A2 => n7, A3 => n61, ZN => p(15));
   U91 : MUX2_X1 port map( A => n12, B => n15, S => A(15), Z => n64);
   U92 : MUX2_X1 port map( A => n10, B => n4, S => A(16), Z => n63);
   U93 : NAND3_X1 port map( A1 => n64, A2 => n7, A3 => n63, ZN => p(16));
   U94 : MUX2_X1 port map( A => n12, B => n15, S => A(16), Z => n66);
   U95 : MUX2_X1 port map( A => n9, B => n4, S => A(17), Z => n65);
   U96 : NAND3_X1 port map( A1 => n66, A2 => n7, A3 => n65, ZN => p(17));
   U97 : MUX2_X1 port map( A => n12, B => n14, S => A(17), Z => n68);
   U98 : MUX2_X1 port map( A => n9, B => n4, S => A(18), Z => n67);
   U99 : NAND3_X1 port map( A1 => n68, A2 => n7, A3 => n67, ZN => p(18));
   U100 : MUX2_X1 port map( A => n12, B => n14, S => A(18), Z => n70);
   U101 : MUX2_X1 port map( A => n9, B => n4, S => A(19), Z => n69);
   U102 : NAND3_X1 port map( A1 => n70, A2 => n7, A3 => n69, ZN => p(19));
   U103 : MUX2_X1 port map( A => n9, B => n4, S => A(20), Z => n71);
   U104 : NAND3_X1 port map( A1 => n72, A2 => n7, A3 => n71, ZN => p(20));
   U105 : MUX2_X1 port map( A => n9, B => n3, S => A(21), Z => n73);
   U106 : NAND3_X1 port map( A1 => n74, A2 => n7, A3 => n73, ZN => p(21));
   U107 : MUX2_X1 port map( A => n9, B => n3, S => A(22), Z => n75);
   U108 : NAND3_X1 port map( A1 => n76, A2 => n7, A3 => n75, ZN => p(22));
   U109 : MUX2_X1 port map( A => n9, B => n3, S => A(23), Z => n77);
   U110 : NAND3_X1 port map( A1 => n78, A2 => n6, A3 => n77, ZN => p(23));
   U111 : MUX2_X1 port map( A => n9, B => n3, S => A(24), Z => n79);
   U112 : NAND3_X1 port map( A1 => n80, A2 => n6, A3 => n79, ZN => p(24));
   U113 : MUX2_X1 port map( A => n14, B => n12, S => n16, Z => n82);
   U114 : MUX2_X1 port map( A => n9, B => n3, S => A(25), Z => n81);
   U115 : NAND3_X1 port map( A1 => n82, A2 => n6, A3 => n81, ZN => p(25));
   U116 : MUX2_X1 port map( A => n14, B => n12, S => n17, Z => n84);
   U117 : MUX2_X1 port map( A => n9, B => n3, S => A(26), Z => n83);
   U118 : NAND3_X1 port map( A1 => n84, A2 => n6, A3 => n83, ZN => p(26));
   U119 : MUX2_X1 port map( A => n14, B => n12, S => n18, Z => n86);
   U120 : MUX2_X1 port map( A => n9, B => n3, S => A(27), Z => n85);
   U121 : NAND3_X1 port map( A1 => n86, A2 => n6, A3 => n85, ZN => p(27));
   U122 : MUX2_X1 port map( A => n14, B => n12, S => n19, Z => n88);
   U123 : MUX2_X1 port map( A => n9, B => n3, S => A(28), Z => n87);
   U124 : NAND3_X1 port map( A1 => n88, A2 => n6, A3 => n87, ZN => p(28));
   U125 : MUX2_X1 port map( A => n14, B => n12, S => n20, Z => n90);
   U126 : MUX2_X1 port map( A => n9, B => n3, S => A(29), Z => n89);
   U127 : NAND3_X1 port map( A1 => n90, A2 => n6, A3 => n89, ZN => p(29));
   U128 : MUX2_X1 port map( A => n14, B => n13, S => n1, Z => n92);
   U129 : MUX2_X1 port map( A => n9, B => n3, S => A(30), Z => n91);
   U130 : NAND3_X1 port map( A1 => n92, A2 => n6, A3 => n91, ZN => p(30));
   U131 : MUX2_X1 port map( A => n14, B => n13, S => n2, Z => n96);
   U132 : MUX2_X1 port map( A => n9, B => n3, S => A(31), Z => n94);
   U133 : NAND3_X1 port map( A1 => n96, A2 => n7, A3 => n94, ZN => p(31));
   U134 : OAI221_X1 port map( B1 => n21, B2 => n14, C1 => A(31), C2 => n11, A 
                           => n9, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_2 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_2;

architecture SYN_beh of ENC_2 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   U3 : BUF_X1 port map( A => n95, Z => n4);
   U4 : BUF_X1 port map( A => n95, Z => n5);
   U5 : BUF_X1 port map( A => n97, Z => n7);
   U6 : BUF_X1 port map( A => n97, Z => n8);
   U7 : BUF_X1 port map( A => n99, Z => n13);
   U8 : BUF_X1 port map( A => n99, Z => n12);
   U9 : BUF_X1 port map( A => n95, Z => n6);
   U10 : BUF_X1 port map( A => n99, Z => n14);
   U11 : MUX2_X1 port map( A => n10, B => n12, S => A(22), Z => n78);
   U12 : BUF_X1 port map( A => n93, Z => n2);
   U13 : BUF_X1 port map( A => n98, Z => n10);
   U14 : MUX2_X1 port map( A => n10, B => n12, S => A(19), Z => n72);
   U15 : MUX2_X1 port map( A => n10, B => n12, S => A(18), Z => n70);
   U16 : MUX2_X1 port map( A => n10, B => n12, S => A(20), Z => n74);
   U17 : MUX2_X1 port map( A => n10, B => n13, S => A(17), Z => n68);
   U18 : MUX2_X1 port map( A => n10, B => n12, S => A(23), Z => n80);
   U19 : BUF_X1 port map( A => n93, Z => n1);
   U20 : BUF_X1 port map( A => n98, Z => n9);
   U21 : MUX2_X1 port map( A => n10, B => n12, S => A(21), Z => n76);
   U22 : BUF_X1 port map( A => n93, Z => n3);
   U23 : BUF_X1 port map( A => n98, Z => n11);
   U24 : INV_X1 port map( A => A(24), ZN => n15);
   U25 : INV_X1 port map( A => A(25), ZN => n16);
   U26 : INV_X1 port map( A => A(26), ZN => n17);
   U27 : INV_X1 port map( A => A(27), ZN => n18);
   U28 : INV_X1 port map( A => A(28), ZN => n19);
   U29 : INV_X1 port map( A => A(29), ZN => n20);
   U30 : INV_X1 port map( A => A(30), ZN => n21);
   U31 : INV_X1 port map( A => A(31), ZN => n22);
   U32 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n27);
   U33 : INV_X1 port map( A => b(2), ZN => n28);
   U34 : INV_X1 port map( A => b(0), ZN => n24);
   U35 : INV_X1 port map( A => b(1), ZN => n23);
   U36 : NAND3_X1 port map( A1 => b(2), A2 => n24, A3 => n23, ZN => n98);
   U37 : NAND2_X1 port map( A1 => b(2), A2 => n27, ZN => n31);
   U38 : XOR2_X1 port map( A => b(1), B => b(0), Z => n25);
   U39 : NAND2_X1 port map( A1 => n25, A2 => n28, ZN => n93);
   U40 : MUX2_X1 port map( A => n31, B => n2, S => A(0), Z => n26);
   U41 : OAI211_X1 port map( C1 => n27, C2 => n28, A => n9, B => n26, ZN => 
                           p(0));
   U42 : INV_X1 port map( A => n27, ZN => n29);
   U43 : NAND2_X1 port map( A1 => n29, A2 => n28, ZN => n99);
   U44 : MUX2_X1 port map( A => n9, B => n13, S => A(0), Z => n34);
   U45 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => n12, ZN => n30);
   U46 : INV_X1 port map( A => n30, ZN => n32);
   U47 : NAND3_X1 port map( A1 => n31, A2 => n1, A3 => n32, ZN => n95);
   U48 : NAND2_X1 port map( A1 => n32, A2 => n1, ZN => n97);
   U49 : MUX2_X1 port map( A => n8, B => n1, S => A(1), Z => n33);
   U50 : NAND3_X1 port map( A1 => n34, A2 => n4, A3 => n33, ZN => p(1));
   U51 : MUX2_X1 port map( A => n9, B => n13, S => A(1), Z => n36);
   U52 : MUX2_X1 port map( A => n8, B => n1, S => A(2), Z => n35);
   U53 : NAND3_X1 port map( A1 => n36, A2 => n6, A3 => n35, ZN => p(2));
   U54 : MUX2_X1 port map( A => n9, B => n13, S => A(2), Z => n38);
   U55 : MUX2_X1 port map( A => n8, B => n1, S => A(3), Z => n37);
   U56 : NAND3_X1 port map( A1 => n38, A2 => n6, A3 => n37, ZN => p(3));
   U57 : MUX2_X1 port map( A => n9, B => n13, S => A(3), Z => n40);
   U58 : MUX2_X1 port map( A => n8, B => n1, S => A(4), Z => n39);
   U59 : NAND3_X1 port map( A1 => n40, A2 => n6, A3 => n39, ZN => p(4));
   U60 : MUX2_X1 port map( A => n9, B => n13, S => A(4), Z => n42);
   U61 : MUX2_X1 port map( A => n8, B => n1, S => A(5), Z => n41);
   U62 : NAND3_X1 port map( A1 => n42, A2 => n6, A3 => n41, ZN => p(5));
   U63 : MUX2_X1 port map( A => n9, B => n13, S => A(5), Z => n44);
   U64 : MUX2_X1 port map( A => n8, B => n1, S => A(6), Z => n43);
   U65 : NAND3_X1 port map( A1 => n44, A2 => n6, A3 => n43, ZN => p(6));
   U66 : MUX2_X1 port map( A => n9, B => n13, S => A(6), Z => n46);
   U67 : MUX2_X1 port map( A => n8, B => n1, S => A(7), Z => n45);
   U68 : NAND3_X1 port map( A1 => n46, A2 => n6, A3 => n45, ZN => p(7));
   U69 : MUX2_X1 port map( A => n9, B => n13, S => A(7), Z => n48);
   U70 : MUX2_X1 port map( A => n8, B => n1, S => A(8), Z => n47);
   U71 : NAND3_X1 port map( A1 => n48, A2 => n5, A3 => n47, ZN => p(8));
   U72 : MUX2_X1 port map( A => n10, B => n13, S => A(8), Z => n50);
   U73 : MUX2_X1 port map( A => n8, B => n1, S => A(9), Z => n49);
   U74 : NAND3_X1 port map( A1 => n50, A2 => n5, A3 => n49, ZN => p(9));
   U75 : MUX2_X1 port map( A => n9, B => n13, S => A(9), Z => n52);
   U76 : MUX2_X1 port map( A => n8, B => n1, S => A(10), Z => n51);
   U77 : NAND3_X1 port map( A1 => n52, A2 => n5, A3 => n51, ZN => p(10));
   U78 : MUX2_X1 port map( A => n9, B => n13, S => A(10), Z => n54);
   U79 : MUX2_X1 port map( A => n8, B => n1, S => A(11), Z => n53);
   U80 : NAND3_X1 port map( A1 => n54, A2 => n5, A3 => n53, ZN => p(11));
   U81 : MUX2_X1 port map( A => n8, B => n1, S => A(12), Z => n56);
   U82 : MUX2_X1 port map( A => n9, B => n13, S => A(11), Z => n55);
   U83 : NAND3_X1 port map( A1 => n6, A2 => n56, A3 => n55, ZN => p(12));
   U84 : MUX2_X1 port map( A => n9, B => n13, S => A(12), Z => n58);
   U85 : MUX2_X1 port map( A => n8, B => n2, S => A(13), Z => n57);
   U86 : NAND3_X1 port map( A1 => n58, A2 => n5, A3 => n57, ZN => p(13));
   U87 : MUX2_X1 port map( A => n9, B => n13, S => A(13), Z => n60);
   U88 : MUX2_X1 port map( A => n8, B => n2, S => A(14), Z => n59);
   U89 : NAND3_X1 port map( A1 => n60, A2 => n5, A3 => n59, ZN => p(14));
   U90 : MUX2_X1 port map( A => n10, B => n14, S => A(14), Z => n62);
   U91 : MUX2_X1 port map( A => n8, B => n2, S => A(15), Z => n61);
   U92 : NAND3_X1 port map( A1 => n62, A2 => n5, A3 => n61, ZN => p(15));
   U93 : MUX2_X1 port map( A => n10, B => n14, S => A(15), Z => n64);
   U94 : MUX2_X1 port map( A => n8, B => n2, S => A(16), Z => n63);
   U95 : NAND3_X1 port map( A1 => n64, A2 => n5, A3 => n63, ZN => p(16));
   U96 : MUX2_X1 port map( A => n10, B => n13, S => A(16), Z => n66);
   U97 : MUX2_X1 port map( A => n7, B => n2, S => A(17), Z => n65);
   U98 : NAND3_X1 port map( A1 => n66, A2 => n5, A3 => n65, ZN => p(17));
   U99 : MUX2_X1 port map( A => n7, B => n2, S => A(18), Z => n67);
   U100 : NAND3_X1 port map( A1 => n68, A2 => n5, A3 => n67, ZN => p(18));
   U101 : MUX2_X1 port map( A => n7, B => n2, S => A(19), Z => n69);
   U102 : NAND3_X1 port map( A1 => n70, A2 => n5, A3 => n69, ZN => p(19));
   U103 : MUX2_X1 port map( A => n7, B => n2, S => A(20), Z => n71);
   U104 : NAND3_X1 port map( A1 => n72, A2 => n4, A3 => n71, ZN => p(20));
   U105 : MUX2_X1 port map( A => n7, B => n2, S => A(21), Z => n73);
   U106 : NAND3_X1 port map( A1 => n74, A2 => n4, A3 => n73, ZN => p(21));
   U107 : MUX2_X1 port map( A => n7, B => n2, S => A(22), Z => n75);
   U108 : NAND3_X1 port map( A1 => n76, A2 => n4, A3 => n75, ZN => p(22));
   U109 : MUX2_X1 port map( A => n7, B => n2, S => A(23), Z => n77);
   U110 : NAND3_X1 port map( A1 => n78, A2 => n4, A3 => n77, ZN => p(23));
   U111 : MUX2_X1 port map( A => n7, B => n2, S => A(24), Z => n79);
   U112 : NAND3_X1 port map( A1 => n80, A2 => n4, A3 => n79, ZN => p(24));
   U113 : MUX2_X1 port map( A => n12, B => n10, S => n15, Z => n82);
   U114 : MUX2_X1 port map( A => n7, B => n2, S => A(25), Z => n81);
   U115 : NAND3_X1 port map( A1 => n82, A2 => n4, A3 => n81, ZN => p(25));
   U116 : MUX2_X1 port map( A => n12, B => n10, S => n16, Z => n84);
   U117 : MUX2_X1 port map( A => n7, B => n2, S => A(26), Z => n83);
   U118 : NAND3_X1 port map( A1 => n84, A2 => n4, A3 => n83, ZN => p(26));
   U119 : MUX2_X1 port map( A => n12, B => n10, S => n17, Z => n86);
   U120 : MUX2_X1 port map( A => n7, B => n2, S => A(27), Z => n85);
   U121 : NAND3_X1 port map( A1 => n86, A2 => n4, A3 => n85, ZN => p(27));
   U122 : MUX2_X1 port map( A => n12, B => n10, S => n18, Z => n88);
   U123 : MUX2_X1 port map( A => n7, B => n3, S => A(28), Z => n87);
   U124 : NAND3_X1 port map( A1 => n88, A2 => n4, A3 => n87, ZN => p(28));
   U125 : MUX2_X1 port map( A => n12, B => n10, S => n19, Z => n90);
   U126 : MUX2_X1 port map( A => n7, B => n3, S => A(29), Z => n89);
   U127 : NAND3_X1 port map( A1 => n90, A2 => n4, A3 => n89, ZN => p(29));
   U128 : MUX2_X1 port map( A => n12, B => n11, S => n20, Z => n92);
   U129 : MUX2_X1 port map( A => n7, B => n3, S => A(30), Z => n91);
   U130 : NAND3_X1 port map( A1 => n92, A2 => n4, A3 => n91, ZN => p(30));
   U131 : MUX2_X1 port map( A => n12, B => n11, S => n21, Z => n96);
   U132 : MUX2_X1 port map( A => n7, B => n1, S => A(31), Z => n94);
   U133 : NAND3_X1 port map( A1 => n96, A2 => n5, A3 => n94, ZN => p(31));
   U134 : OAI221_X1 port map( B1 => n22, B2 => n12, C1 => A(31), C2 => n9, A =>
                           n7, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_1 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_1;

architecture SYN_beh of ENC_1 is

   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96 : std_logic;

begin
   
   U3 : BUF_X1 port map( A => n92, Z => n6);
   U4 : BUF_X1 port map( A => n92, Z => n5);
   U5 : BUF_X1 port map( A => n96, Z => n14);
   U6 : BUF_X1 port map( A => n96, Z => n13);
   U7 : BUF_X1 port map( A => n92, Z => n7);
   U8 : BUF_X1 port map( A => n96, Z => n15);
   U9 : BUF_X1 port map( A => n90, Z => n3);
   U10 : INV_X1 port map( A => n9, ZN => n8);
   U11 : BUF_X1 port map( A => n90, Z => n4);
   U12 : MUX2_X1 port map( A => n11, B => n13, S => A(17), Z => n65);
   U13 : MUX2_X1 port map( A => n11, B => n13, S => A(16), Z => n63);
   U14 : MUX2_X1 port map( A => n11, B => n13, S => A(18), Z => n67);
   U15 : MUX2_X1 port map( A => n11, B => n13, S => A(15), Z => n61);
   U16 : MUX2_X1 port map( A => n11, B => n13, S => A(21), Z => n73);
   U17 : MUX2_X1 port map( A => n11, B => n13, S => A(22), Z => n75);
   U18 : MUX2_X1 port map( A => n11, B => n13, S => A(23), Z => n77);
   U19 : MUX2_X1 port map( A => n11, B => n13, S => A(20), Z => n71);
   U20 : BUF_X1 port map( A => n95, Z => n11);
   U21 : BUF_X1 port map( A => n95, Z => n10);
   U22 : MUX2_X1 port map( A => n11, B => n13, S => A(19), Z => n69);
   U23 : BUF_X1 port map( A => n95, Z => n12);
   U24 : OR2_X1 port map( A1 => b(2), A2 => n24, ZN => n90);
   U25 : XNOR2_X1 port map( A => b(1), B => b(0), ZN => n24);
   U26 : INV_X1 port map( A => A(29), ZN => n1);
   U27 : INV_X1 port map( A => A(30), ZN => n2);
   U28 : INV_X1 port map( A => n94, ZN => n9);
   U29 : INV_X1 port map( A => A(24), ZN => n16);
   U30 : INV_X1 port map( A => A(25), ZN => n17);
   U31 : INV_X1 port map( A => A(26), ZN => n18);
   U32 : INV_X1 port map( A => A(27), ZN => n19);
   U33 : INV_X1 port map( A => A(28), ZN => n20);
   U34 : INV_X1 port map( A => A(31), ZN => n21);
   U35 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n26);
   U36 : INV_X1 port map( A => b(2), ZN => n27);
   U37 : INV_X1 port map( A => b(0), ZN => n23);
   U38 : INV_X1 port map( A => b(1), ZN => n22);
   U39 : NAND3_X1 port map( A1 => b(2), A2 => n23, A3 => n22, ZN => n95);
   U40 : NAND2_X1 port map( A1 => b(2), A2 => n26, ZN => n29);
   U41 : MUX2_X1 port map( A => n29, B => n4, S => A(0), Z => n25);
   U42 : OAI211_X1 port map( C1 => n26, C2 => n27, A => n10, B => n25, ZN => 
                           p(0));
   U43 : INV_X1 port map( A => n26, ZN => n28);
   U44 : NAND2_X1 port map( A1 => n28, A2 => n27, ZN => n96);
   U45 : MUX2_X1 port map( A => n10, B => n14, S => A(0), Z => n31);
   U46 : OAI211_X1 port map( C1 => b(1), C2 => b(0), A => n13, B => n3, ZN => 
                           n94);
   U47 : NAND2_X1 port map( A1 => n9, A2 => n29, ZN => n92);
   U48 : MUX2_X1 port map( A => n94, B => n3, S => A(1), Z => n30);
   U49 : NAND3_X1 port map( A1 => n31, A2 => n5, A3 => n30, ZN => p(1));
   U50 : MUX2_X1 port map( A => n10, B => n15, S => A(1), Z => n33);
   U51 : MUX2_X1 port map( A => n94, B => n3, S => A(2), Z => n32);
   U52 : NAND3_X1 port map( A1 => n33, A2 => n7, A3 => n32, ZN => p(2));
   U53 : MUX2_X1 port map( A => n10, B => n14, S => A(2), Z => n35);
   U54 : MUX2_X1 port map( A => n94, B => n3, S => A(3), Z => n34);
   U55 : NAND3_X1 port map( A1 => n35, A2 => n7, A3 => n34, ZN => p(3));
   U56 : MUX2_X1 port map( A => n10, B => n14, S => A(3), Z => n37);
   U57 : MUX2_X1 port map( A => n94, B => n3, S => A(4), Z => n36);
   U58 : NAND3_X1 port map( A1 => n37, A2 => n7, A3 => n36, ZN => p(4));
   U59 : MUX2_X1 port map( A => n10, B => n14, S => A(4), Z => n39);
   U60 : MUX2_X1 port map( A => n94, B => n3, S => A(5), Z => n38);
   U61 : NAND3_X1 port map( A1 => n39, A2 => n7, A3 => n38, ZN => p(5));
   U62 : MUX2_X1 port map( A => n10, B => n14, S => A(5), Z => n41);
   U63 : MUX2_X1 port map( A => n94, B => n3, S => A(6), Z => n40);
   U64 : NAND3_X1 port map( A1 => n41, A2 => n7, A3 => n40, ZN => p(6));
   U65 : MUX2_X1 port map( A => n10, B => n14, S => A(6), Z => n43);
   U66 : MUX2_X1 port map( A => n94, B => n3, S => A(7), Z => n42);
   U67 : NAND3_X1 port map( A1 => n43, A2 => n7, A3 => n42, ZN => p(7));
   U68 : MUX2_X1 port map( A => n10, B => n14, S => A(7), Z => n45);
   U69 : MUX2_X1 port map( A => n94, B => n3, S => A(8), Z => n44);
   U70 : NAND3_X1 port map( A1 => n45, A2 => n6, A3 => n44, ZN => p(8));
   U71 : MUX2_X1 port map( A => n10, B => n14, S => A(8), Z => n47);
   U72 : MUX2_X1 port map( A => n94, B => n3, S => A(9), Z => n46);
   U73 : NAND3_X1 port map( A1 => n47, A2 => n6, A3 => n46, ZN => p(9));
   U74 : MUX2_X1 port map( A => n94, B => n3, S => A(10), Z => n49);
   U75 : MUX2_X1 port map( A => n10, B => n15, S => A(9), Z => n48);
   U76 : NAND3_X1 port map( A1 => n7, A2 => n49, A3 => n48, ZN => p(10));
   U77 : MUX2_X1 port map( A => n10, B => n14, S => A(10), Z => n51);
   U78 : MUX2_X1 port map( A => n94, B => n3, S => A(11), Z => n50);
   U79 : NAND3_X1 port map( A1 => n51, A2 => n6, A3 => n50, ZN => p(11));
   U80 : MUX2_X1 port map( A => n10, B => n14, S => A(11), Z => n53);
   U81 : MUX2_X1 port map( A => n94, B => n3, S => A(12), Z => n52);
   U82 : NAND3_X1 port map( A1 => n53, A2 => n6, A3 => n52, ZN => p(12));
   U83 : MUX2_X1 port map( A => n10, B => n14, S => A(12), Z => n55);
   U84 : MUX2_X1 port map( A => n94, B => n3, S => A(13), Z => n54);
   U85 : NAND3_X1 port map( A1 => n55, A2 => n6, A3 => n54, ZN => p(13));
   U86 : MUX2_X1 port map( A => n11, B => n14, S => A(13), Z => n57);
   U87 : MUX2_X1 port map( A => n94, B => n3, S => A(14), Z => n56);
   U88 : NAND3_X1 port map( A1 => n57, A2 => n6, A3 => n56, ZN => p(14));
   U89 : MUX2_X1 port map( A => n11, B => n14, S => A(14), Z => n59);
   U90 : MUX2_X1 port map( A => n94, B => n4, S => A(15), Z => n58);
   U91 : NAND3_X1 port map( A1 => n59, A2 => n6, A3 => n58, ZN => p(15));
   U92 : MUX2_X1 port map( A => n8, B => n4, S => A(16), Z => n60);
   U93 : NAND3_X1 port map( A1 => n61, A2 => n6, A3 => n60, ZN => p(16));
   U94 : MUX2_X1 port map( A => n8, B => n4, S => A(17), Z => n62);
   U95 : NAND3_X1 port map( A1 => n63, A2 => n6, A3 => n62, ZN => p(17));
   U96 : MUX2_X1 port map( A => n8, B => n4, S => A(18), Z => n64);
   U97 : NAND3_X1 port map( A1 => n65, A2 => n6, A3 => n64, ZN => p(18));
   U98 : MUX2_X1 port map( A => n8, B => n4, S => A(19), Z => n66);
   U99 : NAND3_X1 port map( A1 => n67, A2 => n6, A3 => n66, ZN => p(19));
   U100 : MUX2_X1 port map( A => n8, B => n4, S => A(20), Z => n68);
   U101 : NAND3_X1 port map( A1 => n69, A2 => n5, A3 => n68, ZN => p(20));
   U102 : MUX2_X1 port map( A => n8, B => n4, S => A(21), Z => n70);
   U103 : NAND3_X1 port map( A1 => n71, A2 => n5, A3 => n70, ZN => p(21));
   U104 : MUX2_X1 port map( A => n8, B => n4, S => A(22), Z => n72);
   U105 : NAND3_X1 port map( A1 => n73, A2 => n5, A3 => n72, ZN => p(22));
   U106 : MUX2_X1 port map( A => n8, B => n4, S => A(23), Z => n74);
   U107 : NAND3_X1 port map( A1 => n75, A2 => n5, A3 => n74, ZN => p(23));
   U108 : MUX2_X1 port map( A => n8, B => n4, S => A(24), Z => n76);
   U109 : NAND3_X1 port map( A1 => n77, A2 => n5, A3 => n76, ZN => p(24));
   U110 : MUX2_X1 port map( A => n13, B => n11, S => n16, Z => n79);
   U111 : MUX2_X1 port map( A => n8, B => n4, S => A(25), Z => n78);
   U112 : NAND3_X1 port map( A1 => n79, A2 => n5, A3 => n78, ZN => p(25));
   U113 : MUX2_X1 port map( A => n13, B => n11, S => n17, Z => n81);
   U114 : MUX2_X1 port map( A => n8, B => n4, S => A(26), Z => n80);
   U115 : NAND3_X1 port map( A1 => n81, A2 => n5, A3 => n80, ZN => p(26));
   U116 : MUX2_X1 port map( A => n14, B => n11, S => n18, Z => n83);
   U117 : MUX2_X1 port map( A => n8, B => n4, S => A(27), Z => n82);
   U118 : NAND3_X1 port map( A1 => n83, A2 => n5, A3 => n82, ZN => p(27));
   U119 : MUX2_X1 port map( A => n14, B => n11, S => n19, Z => n85);
   U120 : MUX2_X1 port map( A => n8, B => n4, S => A(28), Z => n84);
   U121 : NAND3_X1 port map( A1 => n85, A2 => n5, A3 => n84, ZN => p(28));
   U122 : MUX2_X1 port map( A => n14, B => n12, S => n20, Z => n87);
   U123 : MUX2_X1 port map( A => n8, B => n4, S => A(29), Z => n86);
   U124 : NAND3_X1 port map( A1 => n87, A2 => n5, A3 => n86, ZN => p(29));
   U125 : MUX2_X1 port map( A => n13, B => n12, S => n1, Z => n89);
   U126 : MUX2_X1 port map( A => n8, B => n90, S => A(30), Z => n88);
   U127 : NAND3_X1 port map( A1 => n89, A2 => n5, A3 => n88, ZN => p(30));
   U128 : MUX2_X1 port map( A => n13, B => n11, S => n2, Z => n93);
   U129 : MUX2_X1 port map( A => n8, B => n3, S => A(31), Z => n91);
   U130 : NAND3_X1 port map( A1 => n93, A2 => n6, A3 => n91, ZN => p(31));
   U131 : OAI221_X1 port map( B1 => n21, B2 => n13, C1 => A(31), C2 => n10, A 
                           => n8, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPnormalize_SIG_width28_1 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0));

end FPnormalize_SIG_width28_1;

architecture SYN_FPnormalize of FPnormalize_SIG_width28_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n23 : std_logic;

begin
   
   SIG_out(27) <= '0';
   U2 : INV_X2 port map( A => n4, ZN => n2);
   U3 : INV_X2 port map( A => n4, ZN => n3);
   U4 : INV_X1 port map( A => SIG_in(27), ZN => n4);
   U5 : XNOR2_X1 port map( A => EXP_in(6), B => n16, ZN => EXP_out(6));
   U6 : XNOR2_X1 port map( A => EXP_in(7), B => n1, ZN => EXP_out(7));
   U7 : OR2_X1 port map( A1 => n16, A2 => n15, ZN => n1);
   U8 : INV_X1 port map( A => SIG_in(2), ZN => n23);
   U9 : XOR2_X1 port map( A => EXP_in(0), B => n2, Z => EXP_out(0));
   U10 : INV_X1 port map( A => EXP_in(0), ZN => n5);
   U11 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => n6);
   U12 : XOR2_X1 port map( A => EXP_in(1), B => n6, Z => EXP_out(1));
   U13 : NAND3_X1 port map( A1 => EXP_in(1), A2 => n3, A3 => EXP_in(0), ZN => 
                           n7);
   U14 : INV_X1 port map( A => n7, ZN => n10);
   U15 : XOR2_X1 port map( A => EXP_in(2), B => n10, Z => EXP_out(2));
   U16 : INV_X1 port map( A => EXP_in(2), ZN => n8);
   U17 : NOR2_X1 port map( A1 => n8, A2 => n7, ZN => n9);
   U18 : XOR2_X1 port map( A => EXP_in(3), B => n9, Z => EXP_out(3));
   U19 : NAND3_X1 port map( A1 => EXP_in(3), A2 => EXP_in(2), A3 => n10, ZN => 
                           n11);
   U20 : INV_X1 port map( A => n11, ZN => n14);
   U21 : XOR2_X1 port map( A => EXP_in(4), B => n14, Z => EXP_out(4));
   U22 : INV_X1 port map( A => EXP_in(4), ZN => n12);
   U23 : NOR2_X1 port map( A1 => n12, A2 => n11, ZN => n13);
   U24 : XOR2_X1 port map( A => EXP_in(5), B => n13, Z => EXP_out(5));
   U25 : NAND3_X1 port map( A1 => EXP_in(5), A2 => EXP_in(4), A3 => n14, ZN => 
                           n16);
   U26 : INV_X1 port map( A => EXP_in(6), ZN => n15);
   U27 : OAI21_X1 port map( B1 => SIG_in(1), B2 => n4, A => SIG_in(0), ZN => 
                           n17);
   U28 : INV_X1 port map( A => n17, ZN => SIG_out(0));
   U29 : MUX2_X1 port map( A => SIG_in(1), B => SIG_in(2), S => n3, Z => 
                           SIG_out(1));
   U30 : INV_X1 port map( A => SIG_in(3), ZN => n18);
   U31 : MUX2_X1 port map( A => n23, B => n18, S => n3, Z => n19);
   U32 : INV_X1 port map( A => n19, ZN => SIG_out(2));
   U33 : MUX2_X1 port map( A => SIG_in(3), B => SIG_in(4), S => n3, Z => 
                           SIG_out(3));
   U34 : MUX2_X1 port map( A => SIG_in(4), B => SIG_in(5), S => n3, Z => 
                           SIG_out(4));
   U35 : MUX2_X1 port map( A => SIG_in(5), B => SIG_in(6), S => n3, Z => 
                           SIG_out(5));
   U36 : MUX2_X1 port map( A => SIG_in(6), B => SIG_in(7), S => n3, Z => 
                           SIG_out(6));
   U37 : MUX2_X1 port map( A => SIG_in(7), B => SIG_in(8), S => n3, Z => 
                           SIG_out(7));
   U38 : MUX2_X1 port map( A => SIG_in(8), B => SIG_in(9), S => n3, Z => 
                           SIG_out(8));
   U39 : MUX2_X1 port map( A => SIG_in(9), B => SIG_in(10), S => n3, Z => 
                           SIG_out(9));
   U40 : MUX2_X1 port map( A => SIG_in(10), B => SIG_in(11), S => n3, Z => 
                           SIG_out(10));
   U41 : MUX2_X1 port map( A => SIG_in(11), B => SIG_in(12), S => n3, Z => 
                           SIG_out(11));
   U42 : MUX2_X1 port map( A => SIG_in(12), B => SIG_in(13), S => n3, Z => 
                           SIG_out(12));
   U43 : MUX2_X1 port map( A => SIG_in(13), B => SIG_in(14), S => n2, Z => 
                           SIG_out(13));
   U44 : MUX2_X1 port map( A => SIG_in(14), B => SIG_in(15), S => n2, Z => 
                           SIG_out(14));
   U45 : MUX2_X1 port map( A => SIG_in(15), B => SIG_in(16), S => n2, Z => 
                           SIG_out(15));
   U46 : MUX2_X1 port map( A => SIG_in(16), B => SIG_in(17), S => n2, Z => 
                           SIG_out(16));
   U47 : MUX2_X1 port map( A => SIG_in(17), B => SIG_in(18), S => n2, Z => 
                           SIG_out(17));
   U48 : MUX2_X1 port map( A => SIG_in(18), B => SIG_in(19), S => n2, Z => 
                           SIG_out(18));
   U49 : MUX2_X1 port map( A => SIG_in(19), B => SIG_in(20), S => n2, Z => 
                           SIG_out(19));
   U50 : MUX2_X1 port map( A => SIG_in(20), B => SIG_in(21), S => n2, Z => 
                           SIG_out(20));
   U51 : MUX2_X1 port map( A => SIG_in(21), B => SIG_in(22), S => n2, Z => 
                           SIG_out(21));
   U52 : MUX2_X1 port map( A => SIG_in(22), B => SIG_in(23), S => n2, Z => 
                           SIG_out(22));
   U53 : MUX2_X1 port map( A => SIG_in(23), B => SIG_in(24), S => n2, Z => 
                           SIG_out(23));
   U54 : MUX2_X1 port map( A => SIG_in(24), B => SIG_in(25), S => n2, Z => 
                           SIG_out(24));
   U55 : MUX2_X1 port map( A => SIG_in(25), B => SIG_in(26), S => n2, Z => 
                           SIG_out(25));
   U56 : INV_X1 port map( A => SIG_in(26), ZN => n20);
   U57 : NAND2_X1 port map( A1 => n20, A2 => n4, ZN => SIG_out(26));

end SYN_FPnormalize;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity UnpackFP_1 is

   port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector 
         (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, isNaN,
         isINF, isZ, isDN : out std_logic);

end UnpackFP_1;

architecture SYN_UnpackFP of UnpackFP_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, N13, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12
      , n13_port, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37 : std_logic;

begin
   SIG <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, N13, FP(22), 
      FP(21), FP(20), FP(19), FP(18), FP(17), FP(16), FP(15), FP(14), FP(13), 
      FP(12), FP(11), FP(10), FP(9), FP(8), FP(7), FP(6), FP(5), FP(4), FP(3), 
      FP(2), FP(1), FP(0) );
   EXP <= ( FP(30), FP(29), FP(28), FP(27), FP(26), FP(25), FP(24), FP(23) );
   SIGN <= FP(31);
   
   X_Logic0_port <= '0';
   U2 : NAND4_X1 port map( A1 => n24, A2 => n23, A3 => n22, A4 => n21, ZN => 
                           n35);
   U3 : NOR2_X1 port map( A1 => FP(0), A2 => FP(1), ZN => n24);
   U4 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => n22);
   U5 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U6 : NOR2_X1 port map( A1 => FP(10), A2 => FP(9), ZN => n3);
   U7 : INV_X1 port map( A => FP(19), ZN => n17);
   U8 : INV_X1 port map( A => FP(20), ZN => n16);
   U9 : NOR2_X1 port map( A1 => FP(18), A2 => FP(17), ZN => n18);
   U10 : INV_X1 port map( A => FP(13), ZN => n12);
   U11 : INV_X1 port map( A => FP(14), ZN => n11);
   U12 : NOR2_X1 port map( A1 => FP(12), A2 => FP(11), ZN => n13_port);
   U13 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n23);
   U14 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n9);
   U15 : NAND4_X1 port map( A1 => n6, A2 => n5, A3 => n4, A4 => n3, ZN => n10);
   U16 : INV_X1 port map( A => FP(4), ZN => n7);
   U17 : NOR2_X1 port map( A1 => FP(3), A2 => FP(2), ZN => n8);
   U18 : NOR2_X1 port map( A1 => FP(5), A2 => FP(6), ZN => n6);
   U19 : OR2_X1 port map( A1 => FP(22), A2 => FP(21), ZN => n19);
   U20 : OR2_X1 port map( A1 => FP(16), A2 => FP(15), ZN => n14);
   U21 : INV_X1 port map( A => FP(8), ZN => n4);
   U22 : INV_X1 port map( A => FP(7), ZN => n5);
   U23 : NOR4_X1 port map( A1 => FP(27), A2 => FP(28), A3 => FP(29), A4 => 
                           FP(30), ZN => n2);
   U24 : NOR4_X1 port map( A1 => FP(23), A2 => FP(24), A3 => FP(25), A4 => 
                           FP(26), ZN => n1);
   U25 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => N13);
   U26 : NAND3_X1 port map( A1 => n13_port, A2 => n12, A3 => n11, ZN => n15);
   U27 : NAND3_X1 port map( A1 => n18, A2 => n17, A3 => n16, ZN => n20);
   U28 : INV_X1 port map( A => n35, ZN => n37);
   U29 : NOR2_X1 port map( A1 => N13, A2 => n37, ZN => isDN);
   U30 : NOR2_X1 port map( A1 => N13, A2 => n35, ZN => isZ);
   U31 : INV_X1 port map( A => FP(28), ZN => n28);
   U32 : INV_X1 port map( A => FP(27), ZN => n27);
   U33 : INV_X1 port map( A => FP(30), ZN => n26);
   U34 : INV_X1 port map( A => FP(29), ZN => n25);
   U35 : NOR4_X1 port map( A1 => n28, A2 => n27, A3 => n26, A4 => n25, ZN => 
                           n34);
   U36 : INV_X1 port map( A => FP(24), ZN => n32);
   U37 : INV_X1 port map( A => FP(23), ZN => n31);
   U38 : INV_X1 port map( A => FP(26), ZN => n30);
   U39 : INV_X1 port map( A => FP(25), ZN => n29);
   U40 : NOR4_X1 port map( A1 => n32, A2 => n31, A3 => n30, A4 => n29, ZN => 
                           n33);
   U41 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => n36);
   U42 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => isINF);
   U43 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => isNaN);

end SYN_UnpackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_0;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n7, ZN => Y(2));
   U2 : INV_X1 port map( A => n8, ZN => Y(1));
   U3 : INV_X1 port map( A => n9, ZN => Y(0));
   U4 : INV_X1 port map( A => n6, ZN => Y(3));
   U5 : AOI22_X1 port map( A1 => A(2), A2 => SEL, B1 => B(2), B2 => n5, ZN => 
                           n7);
   U6 : AOI22_X1 port map( A1 => A(1), A2 => SEL, B1 => B(1), B2 => n5, ZN => 
                           n8);
   U7 : AOI22_X1 port map( A1 => A(0), A2 => SEL, B1 => B(0), B2 => n5, ZN => 
                           n9);
   U8 : AOI22_X1 port map( A1 => SEL, A2 => A(3), B1 => B(3), B2 => n5, ZN => 
                           n6);
   U9 : INV_X1 port map( A => SEL, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_0;

architecture SYN_STRUCTURAL of RCA_generic_N4_0 is

   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_128 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_127 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_126 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_125 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_0;

architecture SYN_STRUCTURAL of carry_select_N4_0 is

   component MUX21_GENERIC_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1039, n_1040 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1)
                           , A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1039);
   ADDER1 : RCA_generic_N4_31 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1040);
   MUX : MUX21_GENERIC_N4_0 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_0 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_0;

architecture SYN_BEHAVIORAL of PG_GENERAL_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_0 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_0;

architecture SYN_BEHAVIORAL of G_GENERAL_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_0 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_0;

architecture SYN_BEHAVIORAL of PG_NET_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U1 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic_vector 
         (15 downto 0);  S : out std_logic_vector (63 downto 0));

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16;

architecture SYN_STRUCTURAL of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16 is

   component carry_select_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CS_0 : carry_select_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => Ci(0), S(3) => S(3), S(2) 
                           => S(2), S(1) => S(1), S(0) => S(0));
   CS_1 : carry_select_N4_15 port map( A(3) => A(7), A(2) => A(6), A(1) => A(5)
                           , A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1) => 
                           B(5), B(0) => B(4), Ci => Ci(1), S(3) => S(7), S(2) 
                           => S(6), S(1) => S(5), S(0) => S(4));
   CS_2 : carry_select_N4_14 port map( A(3) => A(11), A(2) => A(10), A(1) => 
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Ci => Ci(2), S(3) => 
                           S(11), S(2) => S(10), S(1) => S(9), S(0) => S(8));
   CS_3 : carry_select_N4_13 port map( A(3) => A(15), A(2) => A(14), A(1) => 
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Ci => Ci(3), S(3) => 
                           S(15), S(2) => S(14), S(1) => S(13), S(0) => S(12));
   CS_4 : carry_select_N4_12 port map( A(3) => A(19), A(2) => A(18), A(1) => 
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Ci => Ci(4), S(3) => 
                           S(19), S(2) => S(18), S(1) => S(17), S(0) => S(16));
   CS_5 : carry_select_N4_11 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Ci(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => S(21), S(0) => S(20));
   CS_6 : carry_select_N4_10 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Ci(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CS_7 : carry_select_N4_9 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));
   CS_8 : carry_select_N4_8 port map( A(3) => A(35), A(2) => A(34), A(1) => 
                           A(33), A(0) => A(32), B(3) => B(35), B(2) => B(34), 
                           B(1) => B(33), B(0) => B(32), Ci => Ci(8), S(3) => 
                           S(35), S(2) => S(34), S(1) => S(33), S(0) => S(32));
   CS_9 : carry_select_N4_7 port map( A(3) => A(39), A(2) => A(38), A(1) => 
                           A(37), A(0) => A(36), B(3) => B(39), B(2) => B(38), 
                           B(1) => B(37), B(0) => B(36), Ci => Ci(9), S(3) => 
                           S(39), S(2) => S(38), S(1) => S(37), S(0) => S(36));
   CS_10 : carry_select_N4_6 port map( A(3) => A(43), A(2) => A(42), A(1) => 
                           A(41), A(0) => A(40), B(3) => B(43), B(2) => B(42), 
                           B(1) => B(41), B(0) => B(40), Ci => Ci(10), S(3) => 
                           S(43), S(2) => S(42), S(1) => S(41), S(0) => S(40));
   CS_11 : carry_select_N4_5 port map( A(3) => A(47), A(2) => A(46), A(1) => 
                           A(45), A(0) => A(44), B(3) => B(47), B(2) => B(46), 
                           B(1) => B(45), B(0) => B(44), Ci => Ci(11), S(3) => 
                           S(47), S(2) => S(46), S(1) => S(45), S(0) => S(44));
   CS_12 : carry_select_N4_4 port map( A(3) => A(51), A(2) => A(50), A(1) => 
                           A(49), A(0) => A(48), B(3) => B(51), B(2) => B(50), 
                           B(1) => B(49), B(0) => B(48), Ci => Ci(12), S(3) => 
                           S(51), S(2) => S(50), S(1) => S(49), S(0) => S(48));
   CS_13 : carry_select_N4_3 port map( A(3) => A(55), A(2) => A(54), A(1) => 
                           A(53), A(0) => A(52), B(3) => B(55), B(2) => B(54), 
                           B(1) => B(53), B(0) => B(52), Ci => Ci(13), S(3) => 
                           S(55), S(2) => S(54), S(1) => S(53), S(0) => S(52));
   CS_14 : carry_select_N4_2 port map( A(3) => A(59), A(2) => A(58), A(1) => 
                           A(57), A(0) => A(56), B(3) => B(59), B(2) => B(58), 
                           B(1) => B(57), B(0) => B(56), Ci => Ci(14), S(3) => 
                           S(59), S(2) => S(58), S(1) => S(57), S(0) => S(56));
   CS_15 : carry_select_N4_1 port map( A(3) => A(63), A(2) => A(62), A(1) => 
                           A(61), A(0) => A(60), B(3) => B(63), B(2) => B(62), 
                           B(1) => B(61), B(0) => B(60), Ci => Ci(15), S(3) => 
                           S(63), S(2) => S(62), S(1) => S(61), S(0) => S(60));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (16 downto 0));

end CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_GENERAL_1
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_2
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_3
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_4
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_5
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_6
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_7
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_8
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_1
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_2
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_3
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_4
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_9
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_10
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_11
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_12
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_5
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_6
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_7
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_8
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_9
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_10
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_13
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_14
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_11
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_12
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_13
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_14
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_15
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_16
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_17
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_15
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_18
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_19
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_20
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_21
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_22
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_23
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_24
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_25
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_26
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_27
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_28
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_29
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_30
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_31
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_32
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_16
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_33
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_34
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_35
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_36
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_37
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_38
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_39
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_40
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_41
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_42
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_43
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_44
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_45
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_46
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_47
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_48
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_49
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_50
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_51
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_52
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_53
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_54
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_55
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_56
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_57
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_58
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_59
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_60
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_61
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_62
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_0
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_0
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_NET_1
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_2
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_3
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_4
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_5
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_6
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_7
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_8
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_9
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_10
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_11
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_12
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_13
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_14
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_15
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_16
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_17
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_18
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_19
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_20
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_21
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_22
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_23
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_24
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_25
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_26
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_27
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_28
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_29
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_30
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_31
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_32
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_33
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_34
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_35
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_36
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_37
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_38
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_39
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_40
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_41
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_42
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_43
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_44
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_45
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_46
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_47
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_48
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_49
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_50
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_51
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_52
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_53
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_54
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_55
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_56
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_57
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_58
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_59
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_60
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_61
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_62
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_63
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_0
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   signal Co_16_port, Co_15_port, Co_14_port, Co_13_port, Co_12_port, 
      Co_11_port, Co_10_port, Co_9_port, n8, Co_7_port, Co_6_port, Co_5_port, 
      n9, Co_3_port, Co_2_port, Co_1_port, lev_i_out_5_64_1_port, 
      lev_i_out_5_64_0_port, lev_i_out_5_60_1_port, lev_i_out_5_60_0_port, 
      lev_i_out_5_56_1_port, lev_i_out_5_56_0_port, lev_i_out_5_52_1_port, 
      lev_i_out_5_52_0_port, lev_i_out_4_64_1_port, lev_i_out_4_64_0_port, 
      lev_i_out_4_60_1_port, lev_i_out_4_60_0_port, lev_i_out_4_48_1_port, 
      lev_i_out_4_48_0_port, lev_i_out_4_44_1_port, lev_i_out_4_44_0_port, 
      lev_i_out_4_32_1_port, lev_i_out_4_32_0_port, lev_i_out_4_28_1_port, 
      lev_i_out_4_28_0_port, lev_i_out_3_64_1_port, lev_i_out_3_64_0_port, 
      lev_i_out_3_56_1_port, lev_i_out_3_56_0_port, lev_i_out_3_48_1_port, 
      lev_i_out_3_48_0_port, lev_i_out_3_40_1_port, lev_i_out_3_40_0_port, 
      lev_i_out_3_32_1_port, lev_i_out_3_32_0_port, lev_i_out_3_24_1_port, 
      lev_i_out_3_24_0_port, lev_i_out_3_16_1_port, lev_i_out_3_16_0_port, 
      lev_i_out_2_64_1_port, lev_i_out_2_64_0_port, lev_i_out_2_60_1_port, 
      lev_i_out_2_60_0_port, lev_i_out_2_56_1_port, lev_i_out_2_56_0_port, 
      lev_i_out_2_52_1_port, lev_i_out_2_52_0_port, lev_i_out_2_48_1_port, 
      lev_i_out_2_48_0_port, lev_i_out_2_44_1_port, lev_i_out_2_44_0_port, 
      lev_i_out_2_40_1_port, lev_i_out_2_40_0_port, lev_i_out_2_36_1_port, 
      lev_i_out_2_36_0_port, lev_i_out_2_32_1_port, lev_i_out_2_32_0_port, 
      lev_i_out_2_28_1_port, lev_i_out_2_28_0_port, lev_i_out_2_24_1_port, 
      lev_i_out_2_24_0_port, lev_i_out_2_20_1_port, lev_i_out_2_20_0_port, 
      lev_i_out_2_16_1_port, lev_i_out_2_16_0_port, lev_i_out_2_12_1_port, 
      lev_i_out_2_12_0_port, lev_i_out_2_8_1_port, lev_i_out_2_8_0_port, 
      lev_i_out_1_64_1_port, lev_i_out_1_64_0_port, lev_i_out_1_62_1_port, 
      lev_i_out_1_62_0_port, lev_i_out_1_60_1_port, lev_i_out_1_60_0_port, 
      lev_i_out_1_58_1_port, lev_i_out_1_58_0_port, lev_i_out_1_56_1_port, 
      lev_i_out_1_56_0_port, lev_i_out_1_54_1_port, lev_i_out_1_54_0_port, 
      lev_i_out_1_52_1_port, lev_i_out_1_52_0_port, lev_i_out_1_50_1_port, 
      lev_i_out_1_50_0_port, lev_i_out_1_48_1_port, lev_i_out_1_48_0_port, 
      lev_i_out_1_46_1_port, lev_i_out_1_46_0_port, lev_i_out_1_44_1_port, 
      lev_i_out_1_44_0_port, lev_i_out_1_42_1_port, lev_i_out_1_42_0_port, 
      lev_i_out_1_40_1_port, lev_i_out_1_40_0_port, lev_i_out_1_38_1_port, 
      lev_i_out_1_38_0_port, lev_i_out_1_36_1_port, lev_i_out_1_36_0_port, 
      lev_i_out_1_34_1_port, lev_i_out_1_34_0_port, lev_i_out_1_32_1_port, 
      lev_i_out_1_32_0_port, lev_i_out_1_30_1_port, lev_i_out_1_30_0_port, 
      lev_i_out_1_28_1_port, lev_i_out_1_28_0_port, lev_i_out_1_26_1_port, 
      lev_i_out_1_26_0_port, lev_i_out_1_24_1_port, lev_i_out_1_24_0_port, 
      lev_i_out_1_22_1_port, lev_i_out_1_22_0_port, lev_i_out_1_20_1_port, 
      lev_i_out_1_20_0_port, lev_i_out_1_18_1_port, lev_i_out_1_18_0_port, 
      lev_i_out_1_16_1_port, lev_i_out_1_16_0_port, lev_i_out_1_14_1_port, 
      lev_i_out_1_14_0_port, lev_i_out_1_12_1_port, lev_i_out_1_12_0_port, 
      lev_i_out_1_10_1_port, lev_i_out_1_10_0_port, lev_i_out_1_8_1_port, 
      lev_i_out_1_8_0_port, lev_i_out_1_6_1_port, lev_i_out_1_6_0_port, 
      lev_i_out_1_4_1_port, lev_i_out_1_4_0_port, lev_i_out_1_2_1_port, 
      lev_i_out_0_64_1_port, lev_i_out_0_64_0_port, lev_i_out_0_63_1_port, 
      lev_i_out_0_63_0_port, lev_i_out_0_62_1_port, lev_i_out_0_62_0_port, 
      lev_i_out_0_61_1_port, lev_i_out_0_61_0_port, lev_i_out_0_60_1_port, 
      lev_i_out_0_60_0_port, lev_i_out_0_59_1_port, lev_i_out_0_59_0_port, 
      lev_i_out_0_58_1_port, lev_i_out_0_58_0_port, lev_i_out_0_57_1_port, 
      lev_i_out_0_57_0_port, lev_i_out_0_56_1_port, lev_i_out_0_56_0_port, 
      lev_i_out_0_55_1_port, lev_i_out_0_55_0_port, lev_i_out_0_54_1_port, 
      lev_i_out_0_54_0_port, lev_i_out_0_53_1_port, lev_i_out_0_53_0_port, 
      lev_i_out_0_52_1_port, lev_i_out_0_52_0_port, lev_i_out_0_51_1_port, 
      lev_i_out_0_51_0_port, lev_i_out_0_50_1_port, lev_i_out_0_50_0_port, 
      lev_i_out_0_49_1_port, lev_i_out_0_49_0_port, lev_i_out_0_48_1_port, 
      lev_i_out_0_48_0_port, lev_i_out_0_47_1_port, lev_i_out_0_47_0_port, 
      lev_i_out_0_46_1_port, lev_i_out_0_46_0_port, lev_i_out_0_45_1_port, 
      lev_i_out_0_45_0_port, lev_i_out_0_44_1_port, lev_i_out_0_44_0_port, 
      lev_i_out_0_43_1_port, lev_i_out_0_43_0_port, lev_i_out_0_42_1_port, 
      lev_i_out_0_42_0_port, lev_i_out_0_41_1_port, lev_i_out_0_41_0_port, 
      lev_i_out_0_40_1_port, lev_i_out_0_40_0_port, lev_i_out_0_39_1_port, 
      lev_i_out_0_39_0_port, lev_i_out_0_38_1_port, lev_i_out_0_38_0_port, 
      lev_i_out_0_37_1_port, lev_i_out_0_37_0_port, lev_i_out_0_36_1_port, 
      lev_i_out_0_36_0_port, lev_i_out_0_35_1_port, lev_i_out_0_35_0_port, 
      lev_i_out_0_34_1_port, lev_i_out_0_34_0_port, lev_i_out_0_33_1_port, 
      lev_i_out_0_33_0_port, lev_i_out_0_32_1_port, lev_i_out_0_32_0_port, 
      lev_i_out_0_31_1_port, lev_i_out_0_31_0_port, lev_i_out_0_30_1_port, 
      lev_i_out_0_30_0_port, lev_i_out_0_29_1_port, lev_i_out_0_29_0_port, 
      lev_i_out_0_28_1_port, lev_i_out_0_28_0_port, lev_i_out_0_27_1_port, 
      lev_i_out_0_27_0_port, lev_i_out_0_26_1_port, lev_i_out_0_26_0_port, 
      lev_i_out_0_25_1_port, lev_i_out_0_25_0_port, lev_i_out_0_24_1_port, 
      lev_i_out_0_24_0_port, lev_i_out_0_23_1_port, lev_i_out_0_23_0_port, 
      lev_i_out_0_22_1_port, lev_i_out_0_22_0_port, lev_i_out_0_21_1_port, 
      lev_i_out_0_21_0_port, lev_i_out_0_20_1_port, lev_i_out_0_20_0_port, 
      lev_i_out_0_19_1_port, lev_i_out_0_19_0_port, lev_i_out_0_18_1_port, 
      lev_i_out_0_18_0_port, lev_i_out_0_17_1_port, lev_i_out_0_17_0_port, 
      lev_i_out_0_16_1_port, lev_i_out_0_16_0_port, lev_i_out_0_15_1_port, 
      lev_i_out_0_15_0_port, lev_i_out_0_14_1_port, lev_i_out_0_14_0_port, 
      lev_i_out_0_13_1_port, lev_i_out_0_13_0_port, lev_i_out_0_12_1_port, 
      lev_i_out_0_12_0_port, lev_i_out_0_11_1_port, lev_i_out_0_11_0_port, 
      lev_i_out_0_10_1_port, lev_i_out_0_10_0_port, lev_i_out_0_9_1_port, 
      lev_i_out_0_9_0_port, lev_i_out_0_8_1_port, lev_i_out_0_8_0_port, 
      lev_i_out_0_7_1_port, lev_i_out_0_7_0_port, lev_i_out_0_6_1_port, 
      lev_i_out_0_6_0_port, lev_i_out_0_5_1_port, lev_i_out_0_5_0_port, 
      lev_i_out_0_4_1_port, lev_i_out_0_4_0_port, lev_i_out_0_3_1_port, 
      lev_i_out_0_3_0_port, lev_i_out_0_2_1_port, lev_i_out_0_2_0_port, 
      lev_i_out_0_1_1_port, n1, n2, Co_8_port, Co_4_port, n5, n6, n7, n_1041 : 
      std_logic;

begin
   Co <= ( Co_16_port, Co_15_port, Co_14_port, Co_13_port, Co_12_port, 
      Co_11_port, Co_10_port, Co_9_port, Co_8_port, Co_7_port, Co_6_port, 
      Co_5_port, Co_4_port, Co_3_port, Co_2_port, Co_1_port, Cin );
   
   PG_NETWORK_0_1 : PG_NET_0 port map( A => A(0), B => B(0), G_OUT => 
                           lev_i_out_0_1_1_port, P_OUT => n_1041);
   PG_NETWORK_0_2 : PG_NET_63 port map( A => A(1), B => B(1), G_OUT => 
                           lev_i_out_0_2_1_port, P_OUT => lev_i_out_0_2_0_port)
                           ;
   PG_NETWORK_0_3 : PG_NET_62 port map( A => A(2), B => B(2), G_OUT => 
                           lev_i_out_0_3_1_port, P_OUT => lev_i_out_0_3_0_port)
                           ;
   PG_NETWORK_0_4 : PG_NET_61 port map( A => A(3), B => B(3), G_OUT => 
                           lev_i_out_0_4_1_port, P_OUT => lev_i_out_0_4_0_port)
                           ;
   PG_NETWORK_0_5 : PG_NET_60 port map( A => A(4), B => B(4), G_OUT => 
                           lev_i_out_0_5_1_port, P_OUT => lev_i_out_0_5_0_port)
                           ;
   PG_NETWORK_0_6 : PG_NET_59 port map( A => A(5), B => B(5), G_OUT => 
                           lev_i_out_0_6_1_port, P_OUT => lev_i_out_0_6_0_port)
                           ;
   PG_NETWORK_0_7 : PG_NET_58 port map( A => A(6), B => B(6), G_OUT => 
                           lev_i_out_0_7_1_port, P_OUT => lev_i_out_0_7_0_port)
                           ;
   PG_NETWORK_0_8 : PG_NET_57 port map( A => A(7), B => B(7), G_OUT => 
                           lev_i_out_0_8_1_port, P_OUT => lev_i_out_0_8_0_port)
                           ;
   PG_NETWORK_0_9 : PG_NET_56 port map( A => A(8), B => B(8), G_OUT => 
                           lev_i_out_0_9_1_port, P_OUT => lev_i_out_0_9_0_port)
                           ;
   PG_NETWORK_0_10 : PG_NET_55 port map( A => A(9), B => B(9), G_OUT => 
                           lev_i_out_0_10_1_port, P_OUT => 
                           lev_i_out_0_10_0_port);
   PG_NETWORK_0_11 : PG_NET_54 port map( A => A(10), B => B(10), G_OUT => 
                           lev_i_out_0_11_1_port, P_OUT => 
                           lev_i_out_0_11_0_port);
   PG_NETWORK_0_12 : PG_NET_53 port map( A => A(11), B => B(11), G_OUT => 
                           lev_i_out_0_12_1_port, P_OUT => 
                           lev_i_out_0_12_0_port);
   PG_NETWORK_0_13 : PG_NET_52 port map( A => A(12), B => B(12), G_OUT => 
                           lev_i_out_0_13_1_port, P_OUT => 
                           lev_i_out_0_13_0_port);
   PG_NETWORK_0_14 : PG_NET_51 port map( A => A(13), B => B(13), G_OUT => 
                           lev_i_out_0_14_1_port, P_OUT => 
                           lev_i_out_0_14_0_port);
   PG_NETWORK_0_15 : PG_NET_50 port map( A => A(14), B => B(14), G_OUT => 
                           lev_i_out_0_15_1_port, P_OUT => 
                           lev_i_out_0_15_0_port);
   PG_NETWORK_0_16 : PG_NET_49 port map( A => A(15), B => B(15), G_OUT => 
                           lev_i_out_0_16_1_port, P_OUT => 
                           lev_i_out_0_16_0_port);
   PG_NETWORK_0_17 : PG_NET_48 port map( A => A(16), B => B(16), G_OUT => 
                           lev_i_out_0_17_1_port, P_OUT => 
                           lev_i_out_0_17_0_port);
   PG_NETWORK_0_18 : PG_NET_47 port map( A => A(17), B => B(17), G_OUT => 
                           lev_i_out_0_18_1_port, P_OUT => 
                           lev_i_out_0_18_0_port);
   PG_NETWORK_0_19 : PG_NET_46 port map( A => A(18), B => B(18), G_OUT => 
                           lev_i_out_0_19_1_port, P_OUT => 
                           lev_i_out_0_19_0_port);
   PG_NETWORK_0_20 : PG_NET_45 port map( A => A(19), B => B(19), G_OUT => 
                           lev_i_out_0_20_1_port, P_OUT => 
                           lev_i_out_0_20_0_port);
   PG_NETWORK_0_21 : PG_NET_44 port map( A => A(20), B => B(20), G_OUT => 
                           lev_i_out_0_21_1_port, P_OUT => 
                           lev_i_out_0_21_0_port);
   PG_NETWORK_0_22 : PG_NET_43 port map( A => A(21), B => B(21), G_OUT => 
                           lev_i_out_0_22_1_port, P_OUT => 
                           lev_i_out_0_22_0_port);
   PG_NETWORK_0_23 : PG_NET_42 port map( A => A(22), B => B(22), G_OUT => 
                           lev_i_out_0_23_1_port, P_OUT => 
                           lev_i_out_0_23_0_port);
   PG_NETWORK_0_24 : PG_NET_41 port map( A => A(23), B => B(23), G_OUT => 
                           lev_i_out_0_24_1_port, P_OUT => 
                           lev_i_out_0_24_0_port);
   PG_NETWORK_0_25 : PG_NET_40 port map( A => A(24), B => B(24), G_OUT => 
                           lev_i_out_0_25_1_port, P_OUT => 
                           lev_i_out_0_25_0_port);
   PG_NETWORK_0_26 : PG_NET_39 port map( A => A(25), B => B(25), G_OUT => 
                           lev_i_out_0_26_1_port, P_OUT => 
                           lev_i_out_0_26_0_port);
   PG_NETWORK_0_27 : PG_NET_38 port map( A => A(26), B => B(26), G_OUT => 
                           lev_i_out_0_27_1_port, P_OUT => 
                           lev_i_out_0_27_0_port);
   PG_NETWORK_0_28 : PG_NET_37 port map( A => A(27), B => B(27), G_OUT => 
                           lev_i_out_0_28_1_port, P_OUT => 
                           lev_i_out_0_28_0_port);
   PG_NETWORK_0_29 : PG_NET_36 port map( A => A(28), B => B(28), G_OUT => 
                           lev_i_out_0_29_1_port, P_OUT => 
                           lev_i_out_0_29_0_port);
   PG_NETWORK_0_30 : PG_NET_35 port map( A => A(29), B => B(29), G_OUT => 
                           lev_i_out_0_30_1_port, P_OUT => 
                           lev_i_out_0_30_0_port);
   PG_NETWORK_0_31 : PG_NET_34 port map( A => A(30), B => B(30), G_OUT => 
                           lev_i_out_0_31_1_port, P_OUT => 
                           lev_i_out_0_31_0_port);
   PG_NETWORK_0_32 : PG_NET_33 port map( A => A(31), B => B(31), G_OUT => 
                           lev_i_out_0_32_1_port, P_OUT => 
                           lev_i_out_0_32_0_port);
   PG_NETWORK_0_33 : PG_NET_32 port map( A => A(32), B => B(32), G_OUT => 
                           lev_i_out_0_33_1_port, P_OUT => 
                           lev_i_out_0_33_0_port);
   PG_NETWORK_0_34 : PG_NET_31 port map( A => A(33), B => B(33), G_OUT => 
                           lev_i_out_0_34_1_port, P_OUT => 
                           lev_i_out_0_34_0_port);
   PG_NETWORK_0_35 : PG_NET_30 port map( A => A(34), B => B(34), G_OUT => 
                           lev_i_out_0_35_1_port, P_OUT => 
                           lev_i_out_0_35_0_port);
   PG_NETWORK_0_36 : PG_NET_29 port map( A => A(35), B => B(35), G_OUT => 
                           lev_i_out_0_36_1_port, P_OUT => 
                           lev_i_out_0_36_0_port);
   PG_NETWORK_0_37 : PG_NET_28 port map( A => A(36), B => B(36), G_OUT => 
                           lev_i_out_0_37_1_port, P_OUT => 
                           lev_i_out_0_37_0_port);
   PG_NETWORK_0_38 : PG_NET_27 port map( A => A(37), B => B(37), G_OUT => 
                           lev_i_out_0_38_1_port, P_OUT => 
                           lev_i_out_0_38_0_port);
   PG_NETWORK_0_39 : PG_NET_26 port map( A => A(38), B => B(38), G_OUT => 
                           lev_i_out_0_39_1_port, P_OUT => 
                           lev_i_out_0_39_0_port);
   PG_NETWORK_0_40 : PG_NET_25 port map( A => A(39), B => B(39), G_OUT => 
                           lev_i_out_0_40_1_port, P_OUT => 
                           lev_i_out_0_40_0_port);
   PG_NETWORK_0_41 : PG_NET_24 port map( A => A(40), B => B(40), G_OUT => 
                           lev_i_out_0_41_1_port, P_OUT => 
                           lev_i_out_0_41_0_port);
   PG_NETWORK_0_42 : PG_NET_23 port map( A => A(41), B => B(41), G_OUT => 
                           lev_i_out_0_42_1_port, P_OUT => 
                           lev_i_out_0_42_0_port);
   PG_NETWORK_0_43 : PG_NET_22 port map( A => A(42), B => B(42), G_OUT => 
                           lev_i_out_0_43_1_port, P_OUT => 
                           lev_i_out_0_43_0_port);
   PG_NETWORK_0_44 : PG_NET_21 port map( A => A(43), B => B(43), G_OUT => 
                           lev_i_out_0_44_1_port, P_OUT => 
                           lev_i_out_0_44_0_port);
   PG_NETWORK_0_45 : PG_NET_20 port map( A => A(44), B => B(44), G_OUT => 
                           lev_i_out_0_45_1_port, P_OUT => 
                           lev_i_out_0_45_0_port);
   PG_NETWORK_0_46 : PG_NET_19 port map( A => A(45), B => B(45), G_OUT => 
                           lev_i_out_0_46_1_port, P_OUT => 
                           lev_i_out_0_46_0_port);
   PG_NETWORK_0_47 : PG_NET_18 port map( A => A(46), B => B(46), G_OUT => 
                           lev_i_out_0_47_1_port, P_OUT => 
                           lev_i_out_0_47_0_port);
   PG_NETWORK_0_48 : PG_NET_17 port map( A => A(47), B => B(47), G_OUT => 
                           lev_i_out_0_48_1_port, P_OUT => 
                           lev_i_out_0_48_0_port);
   PG_NETWORK_0_49 : PG_NET_16 port map( A => A(48), B => B(48), G_OUT => 
                           lev_i_out_0_49_1_port, P_OUT => 
                           lev_i_out_0_49_0_port);
   PG_NETWORK_0_50 : PG_NET_15 port map( A => A(49), B => B(49), G_OUT => 
                           lev_i_out_0_50_1_port, P_OUT => 
                           lev_i_out_0_50_0_port);
   PG_NETWORK_0_51 : PG_NET_14 port map( A => A(50), B => B(50), G_OUT => 
                           lev_i_out_0_51_1_port, P_OUT => 
                           lev_i_out_0_51_0_port);
   PG_NETWORK_0_52 : PG_NET_13 port map( A => A(51), B => B(51), G_OUT => 
                           lev_i_out_0_52_1_port, P_OUT => 
                           lev_i_out_0_52_0_port);
   PG_NETWORK_0_53 : PG_NET_12 port map( A => A(52), B => B(52), G_OUT => 
                           lev_i_out_0_53_1_port, P_OUT => 
                           lev_i_out_0_53_0_port);
   PG_NETWORK_0_54 : PG_NET_11 port map( A => A(53), B => B(53), G_OUT => 
                           lev_i_out_0_54_1_port, P_OUT => 
                           lev_i_out_0_54_0_port);
   PG_NETWORK_0_55 : PG_NET_10 port map( A => A(54), B => B(54), G_OUT => 
                           lev_i_out_0_55_1_port, P_OUT => 
                           lev_i_out_0_55_0_port);
   PG_NETWORK_0_56 : PG_NET_9 port map( A => A(55), B => B(55), G_OUT => 
                           lev_i_out_0_56_1_port, P_OUT => 
                           lev_i_out_0_56_0_port);
   PG_NETWORK_0_57 : PG_NET_8 port map( A => A(56), B => B(56), G_OUT => 
                           lev_i_out_0_57_1_port, P_OUT => 
                           lev_i_out_0_57_0_port);
   PG_NETWORK_0_58 : PG_NET_7 port map( A => A(57), B => B(57), G_OUT => 
                           lev_i_out_0_58_1_port, P_OUT => 
                           lev_i_out_0_58_0_port);
   PG_NETWORK_0_59 : PG_NET_6 port map( A => A(58), B => B(58), G_OUT => 
                           lev_i_out_0_59_1_port, P_OUT => 
                           lev_i_out_0_59_0_port);
   PG_NETWORK_0_60 : PG_NET_5 port map( A => A(59), B => B(59), G_OUT => 
                           lev_i_out_0_60_1_port, P_OUT => 
                           lev_i_out_0_60_0_port);
   PG_NETWORK_0_61 : PG_NET_4 port map( A => A(60), B => B(60), G_OUT => 
                           lev_i_out_0_61_1_port, P_OUT => 
                           lev_i_out_0_61_0_port);
   PG_NETWORK_0_62 : PG_NET_3 port map( A => A(61), B => B(61), G_OUT => 
                           lev_i_out_0_62_1_port, P_OUT => 
                           lev_i_out_0_62_0_port);
   PG_NETWORK_0_63 : PG_NET_2 port map( A => A(62), B => B(62), G_OUT => 
                           lev_i_out_0_63_1_port, P_OUT => 
                           lev_i_out_0_63_0_port);
   PG_NETWORK_0_64 : PG_NET_1 port map( A => A(63), B => B(63), G_OUT => 
                           lev_i_out_0_64_1_port, P_OUT => 
                           lev_i_out_0_64_0_port);
   GNET1_1_2 : G_GENERAL_0 port map( PG_ik(1) => lev_i_out_0_2_1_port, PG_ik(0)
                           => lev_i_out_0_2_0_port, G_k_1j => 
                           lev_i_out_0_1_1_port, G_ij => lev_i_out_1_2_1_port);
   PGNET1_1_4 : PG_GENERAL_0 port map( PG_ik(1) => lev_i_out_0_4_1_port, 
                           PG_ik(0) => lev_i_out_0_4_0_port, PG_k_1j(1) => 
                           lev_i_out_0_3_1_port, PG_k_1j(0) => 
                           lev_i_out_0_3_0_port, PG_ij(1) => 
                           lev_i_out_1_4_1_port, PG_ij(0) => 
                           lev_i_out_1_4_0_port);
   PGNET1_1_6 : PG_GENERAL_62 port map( PG_ik(1) => lev_i_out_0_6_1_port, 
                           PG_ik(0) => lev_i_out_0_6_0_port, PG_k_1j(1) => 
                           lev_i_out_0_5_1_port, PG_k_1j(0) => 
                           lev_i_out_0_5_0_port, PG_ij(1) => 
                           lev_i_out_1_6_1_port, PG_ij(0) => 
                           lev_i_out_1_6_0_port);
   PGNET1_1_8 : PG_GENERAL_61 port map( PG_ik(1) => lev_i_out_0_8_1_port, 
                           PG_ik(0) => lev_i_out_0_8_0_port, PG_k_1j(1) => 
                           lev_i_out_0_7_1_port, PG_k_1j(0) => 
                           lev_i_out_0_7_0_port, PG_ij(1) => 
                           lev_i_out_1_8_1_port, PG_ij(0) => 
                           lev_i_out_1_8_0_port);
   PGNET1_1_10 : PG_GENERAL_60 port map( PG_ik(1) => lev_i_out_0_10_1_port, 
                           PG_ik(0) => lev_i_out_0_10_0_port, PG_k_1j(1) => 
                           lev_i_out_0_9_1_port, PG_k_1j(0) => 
                           lev_i_out_0_9_0_port, PG_ij(1) => 
                           lev_i_out_1_10_1_port, PG_ij(0) => 
                           lev_i_out_1_10_0_port);
   PGNET1_1_12 : PG_GENERAL_59 port map( PG_ik(1) => lev_i_out_0_12_1_port, 
                           PG_ik(0) => lev_i_out_0_12_0_port, PG_k_1j(1) => 
                           lev_i_out_0_11_1_port, PG_k_1j(0) => 
                           lev_i_out_0_11_0_port, PG_ij(1) => 
                           lev_i_out_1_12_1_port, PG_ij(0) => 
                           lev_i_out_1_12_0_port);
   PGNET1_1_14 : PG_GENERAL_58 port map( PG_ik(1) => lev_i_out_0_14_1_port, 
                           PG_ik(0) => lev_i_out_0_14_0_port, PG_k_1j(1) => 
                           lev_i_out_0_13_1_port, PG_k_1j(0) => 
                           lev_i_out_0_13_0_port, PG_ij(1) => 
                           lev_i_out_1_14_1_port, PG_ij(0) => 
                           lev_i_out_1_14_0_port);
   PGNET1_1_16 : PG_GENERAL_57 port map( PG_ik(1) => lev_i_out_0_16_1_port, 
                           PG_ik(0) => lev_i_out_0_16_0_port, PG_k_1j(1) => 
                           lev_i_out_0_15_1_port, PG_k_1j(0) => 
                           lev_i_out_0_15_0_port, PG_ij(1) => 
                           lev_i_out_1_16_1_port, PG_ij(0) => 
                           lev_i_out_1_16_0_port);
   PGNET1_1_18 : PG_GENERAL_56 port map( PG_ik(1) => lev_i_out_0_18_1_port, 
                           PG_ik(0) => lev_i_out_0_18_0_port, PG_k_1j(1) => 
                           lev_i_out_0_17_1_port, PG_k_1j(0) => 
                           lev_i_out_0_17_0_port, PG_ij(1) => 
                           lev_i_out_1_18_1_port, PG_ij(0) => 
                           lev_i_out_1_18_0_port);
   PGNET1_1_20 : PG_GENERAL_55 port map( PG_ik(1) => lev_i_out_0_20_1_port, 
                           PG_ik(0) => lev_i_out_0_20_0_port, PG_k_1j(1) => 
                           lev_i_out_0_19_1_port, PG_k_1j(0) => 
                           lev_i_out_0_19_0_port, PG_ij(1) => 
                           lev_i_out_1_20_1_port, PG_ij(0) => 
                           lev_i_out_1_20_0_port);
   PGNET1_1_22 : PG_GENERAL_54 port map( PG_ik(1) => lev_i_out_0_22_1_port, 
                           PG_ik(0) => lev_i_out_0_22_0_port, PG_k_1j(1) => 
                           lev_i_out_0_21_1_port, PG_k_1j(0) => 
                           lev_i_out_0_21_0_port, PG_ij(1) => 
                           lev_i_out_1_22_1_port, PG_ij(0) => 
                           lev_i_out_1_22_0_port);
   PGNET1_1_24 : PG_GENERAL_53 port map( PG_ik(1) => lev_i_out_0_24_1_port, 
                           PG_ik(0) => lev_i_out_0_24_0_port, PG_k_1j(1) => 
                           lev_i_out_0_23_1_port, PG_k_1j(0) => 
                           lev_i_out_0_23_0_port, PG_ij(1) => 
                           lev_i_out_1_24_1_port, PG_ij(0) => 
                           lev_i_out_1_24_0_port);
   PGNET1_1_26 : PG_GENERAL_52 port map( PG_ik(1) => lev_i_out_0_26_1_port, 
                           PG_ik(0) => lev_i_out_0_26_0_port, PG_k_1j(1) => 
                           lev_i_out_0_25_1_port, PG_k_1j(0) => 
                           lev_i_out_0_25_0_port, PG_ij(1) => 
                           lev_i_out_1_26_1_port, PG_ij(0) => 
                           lev_i_out_1_26_0_port);
   PGNET1_1_28 : PG_GENERAL_51 port map( PG_ik(1) => lev_i_out_0_28_1_port, 
                           PG_ik(0) => lev_i_out_0_28_0_port, PG_k_1j(1) => 
                           lev_i_out_0_27_1_port, PG_k_1j(0) => 
                           lev_i_out_0_27_0_port, PG_ij(1) => 
                           lev_i_out_1_28_1_port, PG_ij(0) => 
                           lev_i_out_1_28_0_port);
   PGNET1_1_30 : PG_GENERAL_50 port map( PG_ik(1) => lev_i_out_0_30_1_port, 
                           PG_ik(0) => lev_i_out_0_30_0_port, PG_k_1j(1) => 
                           lev_i_out_0_29_1_port, PG_k_1j(0) => 
                           lev_i_out_0_29_0_port, PG_ij(1) => 
                           lev_i_out_1_30_1_port, PG_ij(0) => 
                           lev_i_out_1_30_0_port);
   PGNET1_1_32 : PG_GENERAL_49 port map( PG_ik(1) => lev_i_out_0_32_1_port, 
                           PG_ik(0) => lev_i_out_0_32_0_port, PG_k_1j(1) => 
                           lev_i_out_0_31_1_port, PG_k_1j(0) => 
                           lev_i_out_0_31_0_port, PG_ij(1) => 
                           lev_i_out_1_32_1_port, PG_ij(0) => 
                           lev_i_out_1_32_0_port);
   PGNET1_1_34 : PG_GENERAL_48 port map( PG_ik(1) => lev_i_out_0_34_1_port, 
                           PG_ik(0) => lev_i_out_0_34_0_port, PG_k_1j(1) => 
                           lev_i_out_0_33_1_port, PG_k_1j(0) => 
                           lev_i_out_0_33_0_port, PG_ij(1) => 
                           lev_i_out_1_34_1_port, PG_ij(0) => 
                           lev_i_out_1_34_0_port);
   PGNET1_1_36 : PG_GENERAL_47 port map( PG_ik(1) => lev_i_out_0_36_1_port, 
                           PG_ik(0) => lev_i_out_0_36_0_port, PG_k_1j(1) => 
                           lev_i_out_0_35_1_port, PG_k_1j(0) => 
                           lev_i_out_0_35_0_port, PG_ij(1) => 
                           lev_i_out_1_36_1_port, PG_ij(0) => 
                           lev_i_out_1_36_0_port);
   PGNET1_1_38 : PG_GENERAL_46 port map( PG_ik(1) => lev_i_out_0_38_1_port, 
                           PG_ik(0) => lev_i_out_0_38_0_port, PG_k_1j(1) => 
                           lev_i_out_0_37_1_port, PG_k_1j(0) => 
                           lev_i_out_0_37_0_port, PG_ij(1) => 
                           lev_i_out_1_38_1_port, PG_ij(0) => 
                           lev_i_out_1_38_0_port);
   PGNET1_1_40 : PG_GENERAL_45 port map( PG_ik(1) => lev_i_out_0_40_1_port, 
                           PG_ik(0) => lev_i_out_0_40_0_port, PG_k_1j(1) => 
                           lev_i_out_0_39_1_port, PG_k_1j(0) => 
                           lev_i_out_0_39_0_port, PG_ij(1) => 
                           lev_i_out_1_40_1_port, PG_ij(0) => 
                           lev_i_out_1_40_0_port);
   PGNET1_1_42 : PG_GENERAL_44 port map( PG_ik(1) => lev_i_out_0_42_1_port, 
                           PG_ik(0) => lev_i_out_0_42_0_port, PG_k_1j(1) => 
                           lev_i_out_0_41_1_port, PG_k_1j(0) => 
                           lev_i_out_0_41_0_port, PG_ij(1) => 
                           lev_i_out_1_42_1_port, PG_ij(0) => 
                           lev_i_out_1_42_0_port);
   PGNET1_1_44 : PG_GENERAL_43 port map( PG_ik(1) => lev_i_out_0_44_1_port, 
                           PG_ik(0) => lev_i_out_0_44_0_port, PG_k_1j(1) => 
                           lev_i_out_0_43_1_port, PG_k_1j(0) => 
                           lev_i_out_0_43_0_port, PG_ij(1) => 
                           lev_i_out_1_44_1_port, PG_ij(0) => 
                           lev_i_out_1_44_0_port);
   PGNET1_1_46 : PG_GENERAL_42 port map( PG_ik(1) => lev_i_out_0_46_1_port, 
                           PG_ik(0) => lev_i_out_0_46_0_port, PG_k_1j(1) => 
                           lev_i_out_0_45_1_port, PG_k_1j(0) => 
                           lev_i_out_0_45_0_port, PG_ij(1) => 
                           lev_i_out_1_46_1_port, PG_ij(0) => 
                           lev_i_out_1_46_0_port);
   PGNET1_1_48 : PG_GENERAL_41 port map( PG_ik(1) => lev_i_out_0_48_1_port, 
                           PG_ik(0) => lev_i_out_0_48_0_port, PG_k_1j(1) => 
                           lev_i_out_0_47_1_port, PG_k_1j(0) => 
                           lev_i_out_0_47_0_port, PG_ij(1) => 
                           lev_i_out_1_48_1_port, PG_ij(0) => 
                           lev_i_out_1_48_0_port);
   PGNET1_1_50 : PG_GENERAL_40 port map( PG_ik(1) => lev_i_out_0_50_1_port, 
                           PG_ik(0) => lev_i_out_0_50_0_port, PG_k_1j(1) => 
                           lev_i_out_0_49_1_port, PG_k_1j(0) => 
                           lev_i_out_0_49_0_port, PG_ij(1) => 
                           lev_i_out_1_50_1_port, PG_ij(0) => 
                           lev_i_out_1_50_0_port);
   PGNET1_1_52 : PG_GENERAL_39 port map( PG_ik(1) => lev_i_out_0_52_1_port, 
                           PG_ik(0) => lev_i_out_0_52_0_port, PG_k_1j(1) => 
                           lev_i_out_0_51_1_port, PG_k_1j(0) => 
                           lev_i_out_0_51_0_port, PG_ij(1) => 
                           lev_i_out_1_52_1_port, PG_ij(0) => 
                           lev_i_out_1_52_0_port);
   PGNET1_1_54 : PG_GENERAL_38 port map( PG_ik(1) => lev_i_out_0_54_1_port, 
                           PG_ik(0) => lev_i_out_0_54_0_port, PG_k_1j(1) => 
                           lev_i_out_0_53_1_port, PG_k_1j(0) => 
                           lev_i_out_0_53_0_port, PG_ij(1) => 
                           lev_i_out_1_54_1_port, PG_ij(0) => 
                           lev_i_out_1_54_0_port);
   PGNET1_1_56 : PG_GENERAL_37 port map( PG_ik(1) => lev_i_out_0_56_1_port, 
                           PG_ik(0) => lev_i_out_0_56_0_port, PG_k_1j(1) => 
                           lev_i_out_0_55_1_port, PG_k_1j(0) => 
                           lev_i_out_0_55_0_port, PG_ij(1) => 
                           lev_i_out_1_56_1_port, PG_ij(0) => 
                           lev_i_out_1_56_0_port);
   PGNET1_1_58 : PG_GENERAL_36 port map( PG_ik(1) => lev_i_out_0_58_1_port, 
                           PG_ik(0) => lev_i_out_0_58_0_port, PG_k_1j(1) => 
                           lev_i_out_0_57_1_port, PG_k_1j(0) => 
                           lev_i_out_0_57_0_port, PG_ij(1) => 
                           lev_i_out_1_58_1_port, PG_ij(0) => 
                           lev_i_out_1_58_0_port);
   PGNET1_1_60 : PG_GENERAL_35 port map( PG_ik(1) => lev_i_out_0_60_1_port, 
                           PG_ik(0) => lev_i_out_0_60_0_port, PG_k_1j(1) => 
                           lev_i_out_0_59_1_port, PG_k_1j(0) => 
                           lev_i_out_0_59_0_port, PG_ij(1) => 
                           lev_i_out_1_60_1_port, PG_ij(0) => 
                           lev_i_out_1_60_0_port);
   PGNET1_1_62 : PG_GENERAL_34 port map( PG_ik(1) => lev_i_out_0_62_1_port, 
                           PG_ik(0) => lev_i_out_0_62_0_port, PG_k_1j(1) => 
                           lev_i_out_0_61_1_port, PG_k_1j(0) => 
                           lev_i_out_0_61_0_port, PG_ij(1) => 
                           lev_i_out_1_62_1_port, PG_ij(0) => 
                           lev_i_out_1_62_0_port);
   PGNET1_1_64 : PG_GENERAL_33 port map( PG_ik(1) => lev_i_out_0_64_1_port, 
                           PG_ik(0) => lev_i_out_0_64_0_port, PG_k_1j(1) => 
                           lev_i_out_0_63_1_port, PG_k_1j(0) => 
                           lev_i_out_0_63_0_port, PG_ij(1) => 
                           lev_i_out_1_64_1_port, PG_ij(0) => 
                           lev_i_out_1_64_0_port);
   GNET_i_2_4_0 : G_GENERAL_16 port map( PG_ik(1) => lev_i_out_1_4_1_port, 
                           PG_ik(0) => lev_i_out_1_4_0_port, G_k_1j => 
                           lev_i_out_1_2_1_port, G_ij => Co_1_port);
   PGNET_i_2_8_0 : PG_GENERAL_32 port map( PG_ik(1) => lev_i_out_1_8_1_port, 
                           PG_ik(0) => lev_i_out_1_8_0_port, PG_k_1j(1) => 
                           lev_i_out_1_6_1_port, PG_k_1j(0) => 
                           lev_i_out_1_6_0_port, PG_ij(1) => 
                           lev_i_out_2_8_1_port, PG_ij(0) => 
                           lev_i_out_2_8_0_port);
   PGNET_i_2_12_0 : PG_GENERAL_31 port map( PG_ik(1) => lev_i_out_1_12_1_port, 
                           PG_ik(0) => lev_i_out_1_12_0_port, PG_k_1j(1) => 
                           lev_i_out_1_10_1_port, PG_k_1j(0) => 
                           lev_i_out_1_10_0_port, PG_ij(1) => 
                           lev_i_out_2_12_1_port, PG_ij(0) => 
                           lev_i_out_2_12_0_port);
   PGNET_i_2_16_0 : PG_GENERAL_30 port map( PG_ik(1) => lev_i_out_1_16_1_port, 
                           PG_ik(0) => lev_i_out_1_16_0_port, PG_k_1j(1) => 
                           lev_i_out_1_14_1_port, PG_k_1j(0) => 
                           lev_i_out_1_14_0_port, PG_ij(1) => 
                           lev_i_out_2_16_1_port, PG_ij(0) => 
                           lev_i_out_2_16_0_port);
   PGNET_i_2_20_0 : PG_GENERAL_29 port map( PG_ik(1) => lev_i_out_1_20_1_port, 
                           PG_ik(0) => lev_i_out_1_20_0_port, PG_k_1j(1) => 
                           lev_i_out_1_18_1_port, PG_k_1j(0) => 
                           lev_i_out_1_18_0_port, PG_ij(1) => 
                           lev_i_out_2_20_1_port, PG_ij(0) => 
                           lev_i_out_2_20_0_port);
   PGNET_i_2_24_0 : PG_GENERAL_28 port map( PG_ik(1) => lev_i_out_1_24_1_port, 
                           PG_ik(0) => lev_i_out_1_24_0_port, PG_k_1j(1) => 
                           lev_i_out_1_22_1_port, PG_k_1j(0) => 
                           lev_i_out_1_22_0_port, PG_ij(1) => 
                           lev_i_out_2_24_1_port, PG_ij(0) => 
                           lev_i_out_2_24_0_port);
   PGNET_i_2_28_0 : PG_GENERAL_27 port map( PG_ik(1) => lev_i_out_1_28_1_port, 
                           PG_ik(0) => lev_i_out_1_28_0_port, PG_k_1j(1) => 
                           lev_i_out_1_26_1_port, PG_k_1j(0) => 
                           lev_i_out_1_26_0_port, PG_ij(1) => 
                           lev_i_out_2_28_1_port, PG_ij(0) => 
                           lev_i_out_2_28_0_port);
   PGNET_i_2_32_0 : PG_GENERAL_26 port map( PG_ik(1) => lev_i_out_1_32_1_port, 
                           PG_ik(0) => lev_i_out_1_32_0_port, PG_k_1j(1) => 
                           lev_i_out_1_30_1_port, PG_k_1j(0) => 
                           lev_i_out_1_30_0_port, PG_ij(1) => 
                           lev_i_out_2_32_1_port, PG_ij(0) => 
                           lev_i_out_2_32_0_port);
   PGNET_i_2_36_0 : PG_GENERAL_25 port map( PG_ik(1) => lev_i_out_1_36_1_port, 
                           PG_ik(0) => lev_i_out_1_36_0_port, PG_k_1j(1) => 
                           lev_i_out_1_34_1_port, PG_k_1j(0) => 
                           lev_i_out_1_34_0_port, PG_ij(1) => 
                           lev_i_out_2_36_1_port, PG_ij(0) => 
                           lev_i_out_2_36_0_port);
   PGNET_i_2_40_0 : PG_GENERAL_24 port map( PG_ik(1) => lev_i_out_1_40_1_port, 
                           PG_ik(0) => lev_i_out_1_40_0_port, PG_k_1j(1) => 
                           lev_i_out_1_38_1_port, PG_k_1j(0) => 
                           lev_i_out_1_38_0_port, PG_ij(1) => 
                           lev_i_out_2_40_1_port, PG_ij(0) => 
                           lev_i_out_2_40_0_port);
   PGNET_i_2_44_0 : PG_GENERAL_23 port map( PG_ik(1) => lev_i_out_1_44_1_port, 
                           PG_ik(0) => lev_i_out_1_44_0_port, PG_k_1j(1) => 
                           lev_i_out_1_42_1_port, PG_k_1j(0) => 
                           lev_i_out_1_42_0_port, PG_ij(1) => 
                           lev_i_out_2_44_1_port, PG_ij(0) => 
                           lev_i_out_2_44_0_port);
   PGNET_i_2_48_0 : PG_GENERAL_22 port map( PG_ik(1) => lev_i_out_1_48_1_port, 
                           PG_ik(0) => lev_i_out_1_48_0_port, PG_k_1j(1) => 
                           lev_i_out_1_46_1_port, PG_k_1j(0) => 
                           lev_i_out_1_46_0_port, PG_ij(1) => 
                           lev_i_out_2_48_1_port, PG_ij(0) => 
                           lev_i_out_2_48_0_port);
   PGNET_i_2_52_0 : PG_GENERAL_21 port map( PG_ik(1) => lev_i_out_1_52_1_port, 
                           PG_ik(0) => lev_i_out_1_52_0_port, PG_k_1j(1) => 
                           lev_i_out_1_50_1_port, PG_k_1j(0) => 
                           lev_i_out_1_50_0_port, PG_ij(1) => 
                           lev_i_out_2_52_1_port, PG_ij(0) => 
                           lev_i_out_2_52_0_port);
   PGNET_i_2_56_0 : PG_GENERAL_20 port map( PG_ik(1) => lev_i_out_1_56_1_port, 
                           PG_ik(0) => lev_i_out_1_56_0_port, PG_k_1j(1) => 
                           lev_i_out_1_54_1_port, PG_k_1j(0) => 
                           lev_i_out_1_54_0_port, PG_ij(1) => 
                           lev_i_out_2_56_1_port, PG_ij(0) => 
                           lev_i_out_2_56_0_port);
   PGNET_i_2_60_0 : PG_GENERAL_19 port map( PG_ik(1) => lev_i_out_1_60_1_port, 
                           PG_ik(0) => lev_i_out_1_60_0_port, PG_k_1j(1) => 
                           lev_i_out_1_58_1_port, PG_k_1j(0) => 
                           lev_i_out_1_58_0_port, PG_ij(1) => 
                           lev_i_out_2_60_1_port, PG_ij(0) => 
                           lev_i_out_2_60_0_port);
   PGNET_i_2_64_0 : PG_GENERAL_18 port map( PG_ik(1) => lev_i_out_1_64_1_port, 
                           PG_ik(0) => lev_i_out_1_64_0_port, PG_k_1j(1) => 
                           lev_i_out_1_62_1_port, PG_k_1j(0) => 
                           lev_i_out_1_62_0_port, PG_ij(1) => 
                           lev_i_out_2_64_1_port, PG_ij(0) => 
                           lev_i_out_2_64_0_port);
   GNET_i_3_8_0 : G_GENERAL_15 port map( PG_ik(1) => lev_i_out_2_8_1_port, 
                           PG_ik(0) => lev_i_out_2_8_0_port, G_k_1j => 
                           Co_1_port, G_ij => Co_2_port);
   PGNET_i_3_16_0 : PG_GENERAL_17 port map( PG_ik(1) => lev_i_out_2_16_1_port, 
                           PG_ik(0) => lev_i_out_2_16_0_port, PG_k_1j(1) => 
                           lev_i_out_2_12_1_port, PG_k_1j(0) => 
                           lev_i_out_2_12_0_port, PG_ij(1) => 
                           lev_i_out_3_16_1_port, PG_ij(0) => 
                           lev_i_out_3_16_0_port);
   PGNET_i_3_24_0 : PG_GENERAL_16 port map( PG_ik(1) => lev_i_out_2_24_1_port, 
                           PG_ik(0) => lev_i_out_2_24_0_port, PG_k_1j(1) => 
                           lev_i_out_2_20_1_port, PG_k_1j(0) => 
                           lev_i_out_2_20_0_port, PG_ij(1) => 
                           lev_i_out_3_24_1_port, PG_ij(0) => 
                           lev_i_out_3_24_0_port);
   PGNET_i_3_32_0 : PG_GENERAL_15 port map( PG_ik(1) => lev_i_out_2_32_1_port, 
                           PG_ik(0) => lev_i_out_2_32_0_port, PG_k_1j(1) => 
                           lev_i_out_2_28_1_port, PG_k_1j(0) => 
                           lev_i_out_2_28_0_port, PG_ij(1) => 
                           lev_i_out_3_32_1_port, PG_ij(0) => 
                           lev_i_out_3_32_0_port);
   PGNET_i_3_40_0 : PG_GENERAL_14 port map( PG_ik(1) => lev_i_out_2_40_1_port, 
                           PG_ik(0) => lev_i_out_2_40_0_port, PG_k_1j(1) => 
                           lev_i_out_2_36_1_port, PG_k_1j(0) => 
                           lev_i_out_2_36_0_port, PG_ij(1) => 
                           lev_i_out_3_40_1_port, PG_ij(0) => 
                           lev_i_out_3_40_0_port);
   PGNET_i_3_48_0 : PG_GENERAL_13 port map( PG_ik(1) => lev_i_out_2_48_1_port, 
                           PG_ik(0) => lev_i_out_2_48_0_port, PG_k_1j(1) => 
                           lev_i_out_2_44_1_port, PG_k_1j(0) => 
                           lev_i_out_2_44_0_port, PG_ij(1) => 
                           lev_i_out_3_48_1_port, PG_ij(0) => 
                           lev_i_out_3_48_0_port);
   PGNET_i_3_56_0 : PG_GENERAL_12 port map( PG_ik(1) => lev_i_out_2_56_1_port, 
                           PG_ik(0) => lev_i_out_2_56_0_port, PG_k_1j(1) => 
                           lev_i_out_2_52_1_port, PG_k_1j(0) => 
                           lev_i_out_2_52_0_port, PG_ij(1) => 
                           lev_i_out_3_56_1_port, PG_ij(0) => 
                           lev_i_out_3_56_0_port);
   PGNET_i_3_64_0 : PG_GENERAL_11 port map( PG_ik(1) => lev_i_out_2_64_1_port, 
                           PG_ik(0) => lev_i_out_2_64_0_port, PG_k_1j(1) => 
                           lev_i_out_2_60_1_port, PG_k_1j(0) => 
                           lev_i_out_2_60_0_port, PG_ij(1) => 
                           lev_i_out_3_64_1_port, PG_ij(0) => 
                           lev_i_out_3_64_0_port);
   GNET_i_4_12_4 : G_GENERAL_14 port map( PG_ik(1) => n1, PG_ik(0) => 
                           lev_i_out_2_12_0_port, G_k_1j => Co_2_port, G_ij => 
                           Co_3_port);
   GNET_i_4_16_0 : G_GENERAL_13 port map( PG_ik(1) => lev_i_out_3_16_1_port, 
                           PG_ik(0) => lev_i_out_3_16_0_port, G_k_1j => 
                           Co_2_port, G_ij => n9);
   PGNET_i_4_28_4 : PG_GENERAL_10 port map( PG_ik(1) => lev_i_out_2_28_1_port, 
                           PG_ik(0) => lev_i_out_2_28_0_port, PG_k_1j(1) => 
                           lev_i_out_3_24_1_port, PG_k_1j(0) => 
                           lev_i_out_3_24_0_port, PG_ij(1) => 
                           lev_i_out_4_28_1_port, PG_ij(0) => 
                           lev_i_out_4_28_0_port);
   PGNET_i_4_32_0 : PG_GENERAL_9 port map( PG_ik(1) => lev_i_out_3_32_1_port, 
                           PG_ik(0) => lev_i_out_3_32_0_port, PG_k_1j(1) => 
                           lev_i_out_3_24_1_port, PG_k_1j(0) => 
                           lev_i_out_3_24_0_port, PG_ij(1) => 
                           lev_i_out_4_32_1_port, PG_ij(0) => 
                           lev_i_out_4_32_0_port);
   PGNET_i_4_44_4 : PG_GENERAL_8 port map( PG_ik(1) => lev_i_out_2_44_1_port, 
                           PG_ik(0) => lev_i_out_2_44_0_port, PG_k_1j(1) => 
                           lev_i_out_3_40_1_port, PG_k_1j(0) => 
                           lev_i_out_3_40_0_port, PG_ij(1) => 
                           lev_i_out_4_44_1_port, PG_ij(0) => 
                           lev_i_out_4_44_0_port);
   PGNET_i_4_48_0 : PG_GENERAL_7 port map( PG_ik(1) => lev_i_out_3_48_1_port, 
                           PG_ik(0) => lev_i_out_3_48_0_port, PG_k_1j(1) => n7,
                           PG_k_1j(0) => lev_i_out_3_40_0_port, PG_ij(1) => 
                           lev_i_out_4_48_1_port, PG_ij(0) => 
                           lev_i_out_4_48_0_port);
   PGNET_i_4_60_4 : PG_GENERAL_6 port map( PG_ik(1) => lev_i_out_2_60_1_port, 
                           PG_ik(0) => lev_i_out_2_60_0_port, PG_k_1j(1) => 
                           lev_i_out_3_56_1_port, PG_k_1j(0) => 
                           lev_i_out_3_56_0_port, PG_ij(1) => 
                           lev_i_out_4_60_1_port, PG_ij(0) => 
                           lev_i_out_4_60_0_port);
   PGNET_i_4_64_0 : PG_GENERAL_5 port map( PG_ik(1) => lev_i_out_3_64_1_port, 
                           PG_ik(0) => lev_i_out_3_64_0_port, PG_k_1j(1) => 
                           lev_i_out_3_56_1_port, PG_k_1j(0) => 
                           lev_i_out_3_56_0_port, PG_ij(1) => 
                           lev_i_out_4_64_1_port, PG_ij(0) => 
                           lev_i_out_4_64_0_port);
   GNET_i_5_20_12 : G_GENERAL_12 port map( PG_ik(1) => lev_i_out_2_20_1_port, 
                           PG_ik(0) => lev_i_out_2_20_0_port, G_k_1j => n9, 
                           G_ij => Co_5_port);
   GNET_i_5_24_8 : G_GENERAL_11 port map( PG_ik(1) => lev_i_out_3_24_1_port, 
                           PG_ik(0) => lev_i_out_3_24_0_port, G_k_1j => n9, 
                           G_ij => Co_6_port);
   GNET_i_5_28_4 : G_GENERAL_10 port map( PG_ik(1) => lev_i_out_4_28_1_port, 
                           PG_ik(0) => lev_i_out_4_28_0_port, G_k_1j => n2, 
                           G_ij => Co_7_port);
   GNET_i_5_32_0 : G_GENERAL_9 port map( PG_ik(1) => lev_i_out_4_32_1_port, 
                           PG_ik(0) => lev_i_out_4_32_0_port, G_k_1j => n9, 
                           G_ij => n8);
   PGNET_i_5_52_12 : PG_GENERAL_4 port map( PG_ik(1) => lev_i_out_2_52_1_port, 
                           PG_ik(0) => lev_i_out_2_52_0_port, PG_k_1j(1) => 
                           lev_i_out_4_48_1_port, PG_k_1j(0) => 
                           lev_i_out_4_48_0_port, PG_ij(1) => 
                           lev_i_out_5_52_1_port, PG_ij(0) => 
                           lev_i_out_5_52_0_port);
   PGNET_i_5_56_8 : PG_GENERAL_3 port map( PG_ik(1) => lev_i_out_3_56_1_port, 
                           PG_ik(0) => lev_i_out_3_56_0_port, PG_k_1j(1) => 
                           lev_i_out_4_48_1_port, PG_k_1j(0) => 
                           lev_i_out_4_48_0_port, PG_ij(1) => 
                           lev_i_out_5_56_1_port, PG_ij(0) => 
                           lev_i_out_5_56_0_port);
   PGNET_i_5_60_4 : PG_GENERAL_2 port map( PG_ik(1) => lev_i_out_4_60_1_port, 
                           PG_ik(0) => lev_i_out_4_60_0_port, PG_k_1j(1) => 
                           lev_i_out_4_48_1_port, PG_k_1j(0) => 
                           lev_i_out_4_48_0_port, PG_ij(1) => 
                           lev_i_out_5_60_1_port, PG_ij(0) => 
                           lev_i_out_5_60_0_port);
   PGNET_i_5_64_0 : PG_GENERAL_1 port map( PG_ik(1) => lev_i_out_4_64_1_port, 
                           PG_ik(0) => lev_i_out_4_64_0_port, PG_k_1j(1) => 
                           lev_i_out_4_48_1_port, PG_k_1j(0) => 
                           lev_i_out_4_48_0_port, PG_ij(1) => 
                           lev_i_out_5_64_1_port, PG_ij(0) => 
                           lev_i_out_5_64_0_port);
   GNET_i_6_36_28 : G_GENERAL_8 port map( PG_ik(1) => n5, PG_ik(0) => 
                           lev_i_out_2_36_0_port, G_k_1j => n8, G_ij => 
                           Co_9_port);
   GNET_i_6_40_24 : G_GENERAL_7 port map( PG_ik(1) => n7, PG_ik(0) => 
                           lev_i_out_3_40_0_port, G_k_1j => n8, G_ij => 
                           Co_10_port);
   GNET_i_6_44_20 : G_GENERAL_6 port map( PG_ik(1) => lev_i_out_4_44_1_port, 
                           PG_ik(0) => lev_i_out_4_44_0_port, G_k_1j => n8, 
                           G_ij => Co_11_port);
   GNET_i_6_48_16 : G_GENERAL_5 port map( PG_ik(1) => lev_i_out_4_48_1_port, 
                           PG_ik(0) => lev_i_out_4_48_0_port, G_k_1j => n6, 
                           G_ij => Co_12_port);
   GNET_i_6_52_12 : G_GENERAL_4 port map( PG_ik(1) => lev_i_out_5_52_1_port, 
                           PG_ik(0) => lev_i_out_5_52_0_port, G_k_1j => n6, 
                           G_ij => Co_13_port);
   GNET_i_6_56_8 : G_GENERAL_3 port map( PG_ik(1) => lev_i_out_5_56_1_port, 
                           PG_ik(0) => lev_i_out_5_56_0_port, G_k_1j => n6, 
                           G_ij => Co_14_port);
   GNET_i_6_60_4 : G_GENERAL_2 port map( PG_ik(1) => lev_i_out_5_60_1_port, 
                           PG_ik(0) => lev_i_out_5_60_0_port, G_k_1j => n6, 
                           G_ij => Co_15_port);
   GNET_i_6_64_0 : G_GENERAL_1 port map( PG_ik(1) => lev_i_out_5_64_1_port, 
                           PG_ik(0) => lev_i_out_5_64_0_port, G_k_1j => n6, 
                           G_ij => Co_16_port);
   U1 : CLKBUF_X1 port map( A => lev_i_out_2_12_1_port, Z => n1);
   U2 : CLKBUF_X1 port map( A => n8, Z => Co_8_port);
   U3 : CLKBUF_X1 port map( A => n9, Z => n2);
   U4 : CLKBUF_X1 port map( A => n2, Z => Co_4_port);
   U5 : CLKBUF_X1 port map( A => lev_i_out_2_36_1_port, Z => n5);
   U6 : CLKBUF_X1 port map( A => Co_8_port, Z => n6);
   U7 : CLKBUF_X1 port map( A => lev_i_out_3_40_1_port, Z => n7);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (63 downto 0);  Cout : out std_logic);

end P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic_vector
            (15 downto 0);  S : out std_logic_vector (63 downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (16 downto 0));
   end component;
   
   signal carry_out_15_port, carry_out_14_port, carry_out_13_port, 
      carry_out_12_port, carry_out_11_port, carry_out_10_port, carry_out_9_port
      , carry_out_8_port, carry_out_7_port, carry_out_6_port, carry_out_5_port,
      carry_out_4_port, carry_out_3_port, carry_out_2_port, carry_out_1_port, 
      carry_out_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38 : std_logic;

begin
   
   CARRY_GEN_INST : CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4 port map( A(63) => 
                           A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => 
                           A(39), A(38) => A(38), A(37) => A(37), A(36) => 
                           A(36), A(35) => A(35), A(34) => A(34), A(33) => 
                           A(33), A(32) => A(32), A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(63) => B(63), B(62) => 
                           B(62), B(61) => B(61), B(60) => B(60), B(59) => 
                           B(59), B(58) => B(58), B(57) => B(57), B(56) => 
                           B(56), B(55) => B(55), B(54) => B(54), B(53) => 
                           B(53), B(52) => B(52), B(51) => B(51), B(50) => 
                           B(50), B(49) => B(49), B(48) => B(48), B(47) => 
                           B(47), B(46) => B(46), B(45) => B(45), B(44) => 
                           B(44), B(43) => B(43), B(42) => B(42), B(41) => 
                           B(41), B(40) => B(40), B(39) => B(39), B(38) => 
                           B(38), B(37) => B(37), B(36) => B(36), B(35) => 
                           B(35), B(34) => B(34), B(33) => B(33), B(32) => 
                           B(32), B(31) => B(31), B(30) => B(30), B(29) => 
                           B(29), B(28) => B(28), B(27) => B(27), B(26) => 
                           B(26), B(25) => B(25), B(24) => B(24), B(23) => 
                           B(23), B(22) => B(22), B(21) => B(21), B(20) => 
                           B(20), B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => B(1), B(0)
                           => B(0), Cin => Cin, Co(16) => Cout, Co(15) => 
                           carry_out_15_port, Co(14) => carry_out_14_port, 
                           Co(13) => carry_out_13_port, Co(12) => 
                           carry_out_12_port, Co(11) => carry_out_11_port, 
                           Co(10) => carry_out_10_port, Co(9) => 
                           carry_out_9_port, Co(8) => carry_out_8_port, Co(7) 
                           => carry_out_7_port, Co(6) => carry_out_6_port, 
                           Co(5) => carry_out_5_port, Co(4) => carry_out_4_port
                           , Co(3) => carry_out_3_port, Co(2) => 
                           carry_out_2_port, Co(1) => carry_out_1_port, Co(0) 
                           => carry_out_0_port);
   SUM_GEN_INST : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16 port map( A(63) => 
                           A(63), A(62) => A(62), A(61) => A(61), A(60) => 
                           A(60), A(59) => A(59), A(58) => A(58), A(57) => 
                           A(57), A(56) => A(56), A(55) => A(55), A(54) => 
                           A(54), A(53) => A(53), A(52) => A(52), A(51) => 
                           A(51), A(50) => A(50), A(49) => A(49), A(48) => 
                           A(48), A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => A(43), A(42) => 
                           A(42), A(41) => A(41), A(40) => A(40), A(39) => n15,
                           A(38) => n19, A(37) => n17, A(36) => n23, A(35) => 
                           n26, A(34) => A(34), A(33) => n16, A(32) => A(32), 
                           A(31) => n38, A(30) => n28, A(29) => n35, A(28) => 
                           A(28), A(27) => n34, A(26) => n18, A(25) => n21, 
                           A(24) => n12, A(23) => n13, A(22) => A(22), A(21) =>
                           n36, A(20) => A(20), A(19) => n8, A(18) => A(18), 
                           A(17) => n37, A(16) => A(16), A(15) => n22, A(14) =>
                           n20, A(13) => n3, A(12) => A(12), A(11) => n1, A(10)
                           => n2, A(9) => A(9), A(8) => A(8), A(7) => A(7), 
                           A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3) => 
                           A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           B(63) => B(63), B(62) => B(62), B(61) => B(61), 
                           B(60) => B(60), B(59) => B(59), B(58) => B(58), 
                           B(57) => B(57), B(56) => B(56), B(55) => B(55), 
                           B(54) => B(54), B(53) => B(53), B(52) => B(52), 
                           B(51) => B(51), B(50) => B(50), B(49) => B(49), 
                           B(48) => B(48), B(47) => B(47), B(46) => B(46), 
                           B(45) => B(45), B(44) => B(44), B(43) => B(43), 
                           B(42) => B(42), B(41) => B(41), B(40) => B(40), 
                           B(39) => n11, B(38) => n9, B(37) => n10, B(36) => 
                           B(36), B(35) => n7, B(34) => B(34), B(33) => n27, 
                           B(32) => B(32), B(31) => n25, B(30) => n32, B(29) =>
                           n24, B(28) => B(28), B(27) => n31, B(26) => n29, 
                           B(25) => n14, B(24) => B(24), B(23) => n33, B(22) =>
                           n6, B(21) => B(21), B(20) => B(20), B(19) => B(19), 
                           B(18) => B(18), B(17) => B(17), B(16) => B(16), 
                           B(15) => n30, B(14) => B(14), B(13) => n5, B(12) => 
                           B(12), B(11) => n4, B(10) => B(10), B(9) => B(9), 
                           B(8) => B(8), B(7) => B(7), B(6) => B(6), B(5) => 
                           B(5), B(4) => B(4), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci(15) => carry_out_15_port, 
                           Ci(14) => carry_out_14_port, Ci(13) => 
                           carry_out_13_port, Ci(12) => carry_out_12_port, 
                           Ci(11) => carry_out_11_port, Ci(10) => 
                           carry_out_10_port, Ci(9) => carry_out_9_port, Ci(8) 
                           => carry_out_8_port, Ci(7) => carry_out_7_port, 
                           Ci(6) => carry_out_6_port, Ci(5) => carry_out_5_port
                           , Ci(4) => carry_out_4_port, Ci(3) => 
                           carry_out_3_port, Ci(2) => carry_out_2_port, Ci(1) 
                           => carry_out_1_port, Ci(0) => carry_out_0_port, 
                           S(63) => S(63), S(62) => S(62), S(61) => S(61), 
                           S(60) => S(60), S(59) => S(59), S(58) => S(58), 
                           S(57) => S(57), S(56) => S(56), S(55) => S(55), 
                           S(54) => S(54), S(53) => S(53), S(52) => S(52), 
                           S(51) => S(51), S(50) => S(50), S(49) => S(49), 
                           S(48) => S(48), S(47) => S(47), S(46) => S(46), 
                           S(45) => S(45), S(44) => S(44), S(43) => S(43), 
                           S(42) => S(42), S(41) => S(41), S(40) => S(40), 
                           S(39) => S(39), S(38) => S(38), S(37) => S(37), 
                           S(36) => S(36), S(35) => S(35), S(34) => S(34), 
                           S(33) => S(33), S(32) => S(32), S(31) => S(31), 
                           S(30) => S(30), S(29) => S(29), S(28) => S(28), 
                           S(27) => S(27), S(26) => S(26), S(25) => S(25), 
                           S(24) => S(24), S(23) => S(23), S(22) => S(22), 
                           S(21) => S(21), S(20) => S(20), S(19) => S(19), 
                           S(18) => S(18), S(17) => S(17), S(16) => S(16), 
                           S(15) => S(15), S(14) => S(14), S(13) => S(13), 
                           S(12) => S(12), S(11) => S(11), S(10) => S(10), S(9)
                           => S(9), S(8) => S(8), S(7) => S(7), S(6) => S(6), 
                           S(5) => S(5), S(4) => S(4), S(3) => S(3), S(2) => 
                           S(2), S(1) => S(1), S(0) => S(0));
   U1 : CLKBUF_X1 port map( A => A(11), Z => n1);
   U2 : CLKBUF_X1 port map( A => A(10), Z => n2);
   U3 : CLKBUF_X1 port map( A => A(13), Z => n3);
   U4 : CLKBUF_X1 port map( A => B(11), Z => n4);
   U5 : CLKBUF_X1 port map( A => B(13), Z => n5);
   U6 : BUF_X1 port map( A => A(24), Z => n12);
   U7 : CLKBUF_X1 port map( A => B(22), Z => n6);
   U8 : CLKBUF_X1 port map( A => B(35), Z => n7);
   U9 : CLKBUF_X1 port map( A => A(19), Z => n8);
   U10 : CLKBUF_X1 port map( A => B(38), Z => n9);
   U11 : CLKBUF_X1 port map( A => A(37), Z => n17);
   U12 : CLKBUF_X1 port map( A => B(37), Z => n10);
   U13 : CLKBUF_X1 port map( A => B(39), Z => n11);
   U14 : BUF_X1 port map( A => B(29), Z => n24);
   U15 : CLKBUF_X1 port map( A => A(23), Z => n13);
   U16 : CLKBUF_X1 port map( A => B(25), Z => n14);
   U17 : CLKBUF_X1 port map( A => A(39), Z => n15);
   U18 : CLKBUF_X1 port map( A => A(33), Z => n16);
   U19 : CLKBUF_X1 port map( A => B(33), Z => n27);
   U20 : CLKBUF_X1 port map( A => A(26), Z => n18);
   U21 : CLKBUF_X1 port map( A => A(38), Z => n19);
   U22 : CLKBUF_X1 port map( A => A(14), Z => n20);
   U23 : CLKBUF_X1 port map( A => A(25), Z => n21);
   U24 : CLKBUF_X1 port map( A => A(15), Z => n22);
   U25 : BUF_X1 port map( A => A(36), Z => n23);
   U26 : CLKBUF_X1 port map( A => B(31), Z => n25);
   U27 : CLKBUF_X1 port map( A => A(35), Z => n26);
   U28 : CLKBUF_X1 port map( A => A(30), Z => n28);
   U29 : CLKBUF_X1 port map( A => A(27), Z => n34);
   U30 : CLKBUF_X1 port map( A => B(26), Z => n29);
   U31 : CLKBUF_X1 port map( A => B(15), Z => n30);
   U32 : CLKBUF_X1 port map( A => B(27), Z => n31);
   U33 : CLKBUF_X1 port map( A => B(30), Z => n32);
   U34 : CLKBUF_X1 port map( A => B(23), Z => n33);
   U35 : CLKBUF_X1 port map( A => A(29), Z => n35);
   U36 : CLKBUF_X1 port map( A => A(21), Z => n36);
   U37 : CLKBUF_X1 port map( A => A(17), Z => n37);
   U38 : CLKBUF_X1 port map( A => A(31), Z => n38);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : INV_X1 port map( A => B, ZN => n4);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U7 : INV_X1 port map( A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_0 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_0;

architecture SYN_rtl of HA_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X2 port map( A1 => B, A2 => A, ZN => C);
   U2 : XOR2_X1 port map( A => A, B => B, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_0 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0));

end ENC_0;

architecture SYN_beh of ENC_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91 : std_logic;

begin
   
   U3 : BUF_X2 port map( A => n86, Z => n11);
   U4 : INV_X1 port map( A => n1, ZN => n51);
   U5 : BUF_X1 port map( A => b(2), Z => n1);
   U6 : BUF_X1 port map( A => b(2), Z => n6);
   U7 : BUF_X4 port map( A => n75, Z => n9);
   U8 : BUF_X1 port map( A => n91, Z => n5);
   U9 : CLKBUF_X3 port map( A => n86, Z => n12);
   U10 : BUF_X1 port map( A => n75, Z => n10);
   U11 : BUF_X2 port map( A => n91, Z => n2);
   U12 : CLKBUF_X1 port map( A => n86, Z => n13);
   U13 : BUF_X1 port map( A => n88, Z => n15);
   U14 : BUF_X1 port map( A => n88, Z => n14);
   U15 : BUF_X1 port map( A => n88, Z => n16);
   U16 : XNOR2_X1 port map( A => n18, B => b(1), ZN => n3);
   U17 : AND2_X1 port map( A1 => n18, A2 => n17, ZN => n4);
   U18 : NAND2_X1 port map( A1 => n3, A2 => n51, ZN => n7);
   U19 : NAND2_X1 port map( A1 => n3, A2 => n51, ZN => n8);
   U20 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n88);
   U21 : INV_X1 port map( A => b(0), ZN => n18);
   U22 : INV_X1 port map( A => b(1), ZN => n17);
   U23 : NAND2_X1 port map( A1 => n4, A2 => n1, ZN => n75);
   U24 : NAND2_X1 port map( A1 => b(2), A2 => n14, ZN => n20);
   U25 : NAND2_X1 port map( A1 => n3, A2 => n51, ZN => n64);
   U26 : MUX2_X1 port map( A => n20, B => n7, S => A(0), Z => n19);
   U27 : OAI211_X1 port map( C1 => n51, C2 => n14, A => n9, B => n19, ZN => 
                           p(0));
   U28 : MUX2_X1 port map( A => n9, B => n14, S => A(0), Z => n22);
   U29 : NAND2_X1 port map( A1 => n6, A2 => n20, ZN => n86);
   U30 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => b(2), ZN => n91);
   U31 : MUX2_X1 port map( A => n5, B => n64, S => A(1), Z => n21);
   U32 : NAND3_X1 port map( A1 => n22, A2 => n11, A3 => n21, ZN => p(1));
   U33 : MUX2_X1 port map( A => n9, B => n14, S => A(1), Z => n24);
   U34 : MUX2_X1 port map( A => n2, B => n8, S => A(2), Z => n23);
   U35 : NAND3_X1 port map( A1 => n24, A2 => n13, A3 => n23, ZN => p(2));
   U36 : MUX2_X1 port map( A => n9, B => n14, S => A(2), Z => n26);
   U37 : MUX2_X1 port map( A => n2, B => n84, S => A(3), Z => n25);
   U38 : NAND3_X1 port map( A1 => n26, A2 => n13, A3 => n25, ZN => p(3));
   U39 : MUX2_X1 port map( A => n9, B => n14, S => A(3), Z => n28);
   U40 : MUX2_X1 port map( A => n5, B => n7, S => A(4), Z => n27);
   U41 : NAND3_X1 port map( A1 => n28, A2 => n13, A3 => n27, ZN => p(4));
   U42 : MUX2_X1 port map( A => n9, B => n14, S => A(4), Z => n30);
   U43 : MUX2_X1 port map( A => n2, B => n64, S => A(5), Z => n29);
   U44 : NAND3_X1 port map( A1 => n30, A2 => n13, A3 => n29, ZN => p(5));
   U45 : MUX2_X1 port map( A => n9, B => n14, S => A(5), Z => n32);
   U46 : MUX2_X1 port map( A => n2, B => n8, S => A(6), Z => n31);
   U47 : NAND3_X1 port map( A1 => n32, A2 => n13, A3 => n31, ZN => p(6));
   U48 : MUX2_X1 port map( A => n9, B => n14, S => A(6), Z => n34);
   U49 : MUX2_X1 port map( A => n5, B => n84, S => A(7), Z => n33);
   U50 : NAND3_X1 port map( A1 => n34, A2 => n13, A3 => n33, ZN => p(7));
   U51 : MUX2_X1 port map( A => n9, B => n14, S => A(7), Z => n36);
   U52 : MUX2_X1 port map( A => n2, B => n8, S => A(8), Z => n35);
   U53 : NAND3_X1 port map( A1 => n36, A2 => n12, A3 => n35, ZN => p(8));
   U54 : MUX2_X1 port map( A => n9, B => n14, S => A(8), Z => n38);
   U55 : MUX2_X1 port map( A => n5, B => n64, S => A(9), Z => n37);
   U56 : NAND3_X1 port map( A1 => n38, A2 => n12, A3 => n37, ZN => p(9));
   U57 : MUX2_X1 port map( A => n9, B => n14, S => A(9), Z => n40);
   U58 : MUX2_X1 port map( A => n2, B => n7, S => A(10), Z => n39);
   U59 : NAND3_X1 port map( A1 => n40, A2 => n12, A3 => n39, ZN => p(10));
   U60 : MUX2_X1 port map( A => n9, B => n14, S => A(10), Z => n42);
   U61 : MUX2_X1 port map( A => n2, B => n7, S => A(11), Z => n41);
   U62 : NAND3_X1 port map( A1 => n42, A2 => n12, A3 => n41, ZN => p(11));
   U63 : MUX2_X1 port map( A => n9, B => n14, S => A(11), Z => n44);
   U64 : MUX2_X1 port map( A => n2, B => n8, S => A(12), Z => n43);
   U65 : NAND3_X1 port map( A1 => n44, A2 => n12, A3 => n43, ZN => p(12));
   U66 : MUX2_X1 port map( A => n9, B => n14, S => A(12), Z => n46);
   U67 : MUX2_X1 port map( A => n5, B => n64, S => A(13), Z => n45);
   U68 : NAND3_X1 port map( A1 => n46, A2 => n12, A3 => n45, ZN => p(13));
   U69 : MUX2_X1 port map( A => n9, B => n15, S => A(13), Z => n48);
   U70 : MUX2_X1 port map( A => n2, B => n84, S => A(14), Z => n47);
   U71 : NAND3_X1 port map( A1 => n48, A2 => n12, A3 => n47, ZN => p(14));
   U72 : MUX2_X1 port map( A => n2, B => n84, S => A(15), Z => n50);
   U73 : MUX2_X1 port map( A => n9, B => n15, S => A(14), Z => n49);
   U74 : NAND3_X1 port map( A1 => n13, A2 => n50, A3 => n49, ZN => p(15));
   U75 : MUX2_X1 port map( A => n9, B => n15, S => A(15), Z => n53);
   U76 : NAND2_X1 port map( A1 => n3, A2 => n51, ZN => n84);
   U77 : MUX2_X1 port map( A => n2, B => n84, S => A(16), Z => n52);
   U78 : NAND3_X1 port map( A1 => n53, A2 => n12, A3 => n52, ZN => p(16));
   U79 : MUX2_X1 port map( A => n9, B => n15, S => A(16), Z => n55);
   U80 : MUX2_X1 port map( A => n2, B => n7, S => A(17), Z => n54);
   U81 : NAND3_X1 port map( A1 => n55, A2 => n12, A3 => n54, ZN => p(17));
   U82 : MUX2_X1 port map( A => n9, B => n15, S => A(17), Z => n57);
   U83 : MUX2_X1 port map( A => n2, B => n64, S => A(18), Z => n56);
   U84 : NAND3_X1 port map( A1 => n57, A2 => n12, A3 => n56, ZN => p(18));
   U85 : MUX2_X1 port map( A => n9, B => n15, S => A(18), Z => n59);
   U86 : MUX2_X1 port map( A => n5, B => n8, S => A(19), Z => n58);
   U87 : NAND3_X1 port map( A1 => n59, A2 => n12, A3 => n58, ZN => p(19));
   U88 : MUX2_X1 port map( A => n9, B => n15, S => A(19), Z => n61);
   U89 : MUX2_X1 port map( A => n2, B => n8, S => A(20), Z => n60);
   U90 : NAND3_X1 port map( A1 => n61, A2 => n11, A3 => n60, ZN => p(20));
   U91 : MUX2_X1 port map( A => n9, B => n15, S => A(20), Z => n63);
   U92 : MUX2_X1 port map( A => n2, B => n64, S => A(21), Z => n62);
   U93 : NAND3_X1 port map( A1 => n63, A2 => n11, A3 => n62, ZN => p(21));
   U94 : MUX2_X1 port map( A => n9, B => n15, S => A(21), Z => n66);
   U95 : MUX2_X1 port map( A => n2, B => n7, S => A(22), Z => n65);
   U96 : NAND3_X1 port map( A1 => n66, A2 => n11, A3 => n65, ZN => p(22));
   U97 : MUX2_X1 port map( A => n5, B => n64, S => A(23), Z => n68);
   U98 : MUX2_X1 port map( A => n10, B => n15, S => A(22), Z => n67);
   U99 : NAND3_X1 port map( A1 => n68, A2 => n11, A3 => n67, ZN => p(23));
   U100 : MUX2_X1 port map( A => n10, B => n15, S => A(23), Z => n70);
   U101 : MUX2_X1 port map( A => n2, B => n7, S => A(24), Z => n69);
   U102 : NAND3_X1 port map( A1 => n70, A2 => n11, A3 => n69, ZN => p(24));
   U103 : MUX2_X1 port map( A => n10, B => n15, S => A(24), Z => n72);
   U104 : MUX2_X1 port map( A => n2, B => n84, S => A(25), Z => n71);
   U105 : NAND3_X1 port map( A1 => n72, A2 => n11, A3 => n71, ZN => p(25));
   U106 : MUX2_X1 port map( A => n2, B => n8, S => A(26), Z => n74);
   U107 : NAND2_X1 port map( A1 => n4, A2 => n6, ZN => n89);
   U108 : MUX2_X1 port map( A => n89, B => n15, S => A(25), Z => n73);
   U109 : NAND3_X1 port map( A1 => n74, A2 => n73, A3 => n11, ZN => p(26));
   U110 : MUX2_X1 port map( A => n10, B => n15, S => A(26), Z => n77);
   U111 : MUX2_X1 port map( A => n2, B => n64, S => A(27), Z => n76);
   U112 : NAND3_X1 port map( A1 => n77, A2 => n11, A3 => n76, ZN => p(27));
   U113 : MUX2_X1 port map( A => n89, B => n15, S => A(27), Z => n79);
   U114 : MUX2_X1 port map( A => n5, B => n7, S => A(28), Z => n78);
   U115 : NAND3_X1 port map( A1 => n79, A2 => n11, A3 => n78, ZN => p(28));
   U116 : MUX2_X1 port map( A => n89, B => n15, S => A(28), Z => n81);
   U117 : MUX2_X1 port map( A => n91, B => n84, S => A(29), Z => n80);
   U118 : NAND3_X1 port map( A1 => n81, A2 => n11, A3 => n80, ZN => p(29));
   U119 : MUX2_X1 port map( A => n10, B => n16, S => A(29), Z => n83);
   U120 : MUX2_X1 port map( A => n5, B => n84, S => A(30), Z => n82);
   U121 : NAND3_X1 port map( A1 => n83, A2 => n11, A3 => n82, ZN => p(30));
   U122 : MUX2_X1 port map( A => n89, B => n16, S => A(30), Z => n87);
   U123 : MUX2_X1 port map( A => n5, B => n8, S => A(31), Z => n85);
   U124 : NAND3_X1 port map( A1 => n85, A2 => n12, A3 => n87, ZN => p(31));
   U125 : MUX2_X1 port map( A => n89, B => n16, S => A(31), Z => n90);
   U126 : NAND2_X1 port map( A1 => n5, A2 => n90, ZN => p(32));

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PackFP is

   port( SIGN : in std_logic;  EXP : in std_logic_vector (7 downto 0);  SIG : 
         in std_logic_vector (22 downto 0);  isNaN, isINF, isZ : in std_logic; 
         FP : out std_logic_vector (31 downto 0));

end PackFP;

architecture SYN_PackFP of PackFP is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal FP_30_port, FP_29_port, FP_28_port, FP_27_port, FP_26_port, 
      FP_25_port, FP_24_port, FP_23_port, FP_22_port, FP_21_port, FP_20_port, 
      FP_19_port, FP_18_port, FP_17_port, FP_16_port, FP_15_port, FP_14_port, 
      FP_13_port, FP_12_port, FP_11_port, FP_10_port, FP_9_port, FP_8_port, 
      FP_7_port, FP_6_port, FP_5_port, FP_4_port, FP_3_port, FP_2_port, 
      FP_1_port, FP_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15 : std_logic;

begin
   FP <= ( SIGN, FP_30_port, FP_29_port, FP_28_port, FP_27_port, FP_26_port, 
      FP_25_port, FP_24_port, FP_23_port, FP_22_port, FP_21_port, FP_20_port, 
      FP_19_port, FP_18_port, FP_17_port, FP_16_port, FP_15_port, FP_14_port, 
      FP_13_port, FP_12_port, FP_11_port, FP_10_port, FP_9_port, FP_8_port, 
      FP_7_port, FP_6_port, FP_5_port, FP_4_port, FP_3_port, FP_2_port, 
      FP_1_port, FP_0_port );
   
   U3 : AND2_X2 port map( A1 => n2, A2 => n14, ZN => n1);
   U4 : NAND2_X2 port map( A1 => n3, A2 => n5, ZN => n13);
   U5 : INV_X2 port map( A => isZ, ZN => n14);
   U6 : INV_X1 port map( A => isINF, ZN => n3);
   U7 : INV_X1 port map( A => isNaN, ZN => n5);
   U8 : INV_X1 port map( A => n13, ZN => n2);
   U9 : AND2_X1 port map( A1 => SIG(0), A2 => n1, ZN => FP_0_port);
   U10 : AND2_X1 port map( A1 => SIG(1), A2 => n1, ZN => FP_1_port);
   U11 : AND2_X1 port map( A1 => SIG(2), A2 => n1, ZN => FP_2_port);
   U12 : AND2_X1 port map( A1 => SIG(3), A2 => n1, ZN => FP_3_port);
   U13 : AND2_X1 port map( A1 => SIG(4), A2 => n1, ZN => FP_4_port);
   U14 : AND2_X1 port map( A1 => SIG(5), A2 => n1, ZN => FP_5_port);
   U15 : AND2_X1 port map( A1 => SIG(6), A2 => n1, ZN => FP_6_port);
   U16 : AND2_X1 port map( A1 => SIG(7), A2 => n1, ZN => FP_7_port);
   U17 : AND2_X1 port map( A1 => SIG(8), A2 => n1, ZN => FP_8_port);
   U18 : AND2_X1 port map( A1 => SIG(9), A2 => n1, ZN => FP_9_port);
   U19 : AND2_X1 port map( A1 => SIG(10), A2 => n1, ZN => FP_10_port);
   U20 : AND2_X1 port map( A1 => SIG(11), A2 => n1, ZN => FP_11_port);
   U21 : AND2_X1 port map( A1 => SIG(12), A2 => n1, ZN => FP_12_port);
   U22 : AND2_X1 port map( A1 => SIG(13), A2 => n1, ZN => FP_13_port);
   U23 : AND2_X1 port map( A1 => SIG(14), A2 => n1, ZN => FP_14_port);
   U24 : AND2_X1 port map( A1 => SIG(15), A2 => n1, ZN => FP_15_port);
   U25 : AND2_X1 port map( A1 => SIG(16), A2 => n1, ZN => FP_16_port);
   U26 : AND2_X1 port map( A1 => SIG(17), A2 => n1, ZN => FP_17_port);
   U27 : AND2_X1 port map( A1 => SIG(18), A2 => n1, ZN => FP_18_port);
   U28 : AND2_X1 port map( A1 => SIG(19), A2 => n1, ZN => FP_19_port);
   U29 : AND2_X1 port map( A1 => SIG(20), A2 => n1, ZN => FP_20_port);
   U30 : AND2_X1 port map( A1 => SIG(21), A2 => n1, ZN => FP_21_port);
   U31 : NAND3_X1 port map( A1 => SIG(22), A2 => n3, A3 => n14, ZN => n4);
   U32 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => FP_22_port);
   U33 : AOI21_X1 port map( B1 => EXP(0), B2 => n14, A => n13, ZN => n6);
   U34 : INV_X1 port map( A => n6, ZN => FP_23_port);
   U35 : AOI21_X1 port map( B1 => EXP(1), B2 => n14, A => n13, ZN => n7);
   U36 : INV_X1 port map( A => n7, ZN => FP_24_port);
   U37 : AOI21_X1 port map( B1 => EXP(2), B2 => n14, A => n13, ZN => n8);
   U38 : INV_X1 port map( A => n8, ZN => FP_25_port);
   U39 : AOI21_X1 port map( B1 => EXP(3), B2 => n14, A => n13, ZN => n9);
   U40 : INV_X1 port map( A => n9, ZN => FP_26_port);
   U41 : AOI21_X1 port map( B1 => EXP(4), B2 => n14, A => n13, ZN => n10);
   U42 : INV_X1 port map( A => n10, ZN => FP_27_port);
   U43 : AOI21_X1 port map( B1 => EXP(5), B2 => n14, A => n13, ZN => n11);
   U44 : INV_X1 port map( A => n11, ZN => FP_28_port);
   U45 : AOI21_X1 port map( B1 => EXP(6), B2 => n14, A => n13, ZN => n12);
   U46 : INV_X1 port map( A => n12, ZN => FP_29_port);
   U47 : AOI21_X1 port map( B1 => EXP(7), B2 => n14, A => n13, ZN => n15);
   U48 : INV_X1 port map( A => n15, ZN => FP_30_port);

end SYN_PackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPround_SIG_width28 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0));

end FPround_SIG_width28;

architecture SYN_FPround of FPround_SIG_width28 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FPround_SIG_width28_DW01_inc_1
      port( A : in std_logic_vector (24 downto 0);  SUM : out std_logic_vector 
            (24 downto 0));
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, n1, n2_port, n3_port : 
      std_logic;

begin
   EXP_out <= ( EXP_in(7), EXP_in(6), EXP_in(5), EXP_in(4), EXP_in(3), 
      EXP_in(2), EXP_in(1), EXP_in(0) );
   
   SIG_out(2) <= '0';
   add_45 : FPround_SIG_width28_DW01_inc_1 port map( A(24) => SIG_in(27), A(23)
                           => SIG_in(26), A(22) => SIG_in(25), A(21) => 
                           SIG_in(24), A(20) => SIG_in(23), A(19) => SIG_in(22)
                           , A(18) => SIG_in(21), A(17) => SIG_in(20), A(16) =>
                           SIG_in(19), A(15) => SIG_in(18), A(14) => SIG_in(17)
                           , A(13) => SIG_in(16), A(12) => SIG_in(15), A(11) =>
                           SIG_in(14), A(10) => SIG_in(13), A(9) => SIG_in(12),
                           A(8) => SIG_in(11), A(7) => SIG_in(10), A(6) => 
                           SIG_in(9), A(5) => SIG_in(8), A(4) => SIG_in(7), 
                           A(3) => SIG_in(6), A(2) => SIG_in(5), A(1) => 
                           SIG_in(4), A(0) => SIG_in(3), SUM(24) => N26, 
                           SUM(23) => N25, SUM(22) => N24, SUM(21) => N23, 
                           SUM(20) => N22, SUM(19) => N21, SUM(18) => N20, 
                           SUM(17) => N19, SUM(16) => N18, SUM(15) => N17, 
                           SUM(14) => N16, SUM(13) => N15, SUM(12) => N14, 
                           SUM(11) => N13, SUM(10) => N12, SUM(9) => N11, 
                           SUM(8) => N10, SUM(7) => N9, SUM(6) => N8, SUM(5) =>
                           N7, SUM(4) => N6, SUM(3) => N5, SUM(2) => N4, SUM(1)
                           => N3, SUM(0) => N2);
   U3 : INV_X1 port map( A => n3_port, ZN => n1);
   U4 : INV_X1 port map( A => n3_port, ZN => n2_port);
   U5 : INV_X1 port map( A => SIG_in(2), ZN => n3_port);
   U6 : AND2_X1 port map( A1 => SIG_in(0), A2 => n3_port, ZN => SIG_out(0));
   U7 : AND2_X1 port map( A1 => SIG_in(1), A2 => n3_port, ZN => SIG_out(1));
   U8 : MUX2_X1 port map( A => SIG_in(3), B => N2, S => n1, Z => SIG_out(3));
   U9 : MUX2_X1 port map( A => SIG_in(4), B => N3, S => n1, Z => SIG_out(4));
   U10 : MUX2_X1 port map( A => SIG_in(5), B => N4, S => n1, Z => SIG_out(5));
   U11 : MUX2_X1 port map( A => SIG_in(6), B => N5, S => n1, Z => SIG_out(6));
   U12 : MUX2_X1 port map( A => SIG_in(7), B => N6, S => n1, Z => SIG_out(7));
   U13 : MUX2_X1 port map( A => SIG_in(8), B => N7, S => n1, Z => SIG_out(8));
   U14 : MUX2_X1 port map( A => SIG_in(9), B => N8, S => n1, Z => SIG_out(9));
   U15 : MUX2_X1 port map( A => SIG_in(10), B => N9, S => n1, Z => SIG_out(10))
                           ;
   U16 : MUX2_X1 port map( A => SIG_in(11), B => N10, S => n1, Z => SIG_out(11)
                           );
   U17 : MUX2_X1 port map( A => SIG_in(12), B => N11, S => n1, Z => SIG_out(12)
                           );
   U18 : MUX2_X1 port map( A => SIG_in(13), B => N12, S => n1, Z => SIG_out(13)
                           );
   U19 : MUX2_X1 port map( A => SIG_in(14), B => N13, S => n1, Z => SIG_out(14)
                           );
   U20 : MUX2_X1 port map( A => SIG_in(15), B => N14, S => n2_port, Z => 
                           SIG_out(15));
   U21 : MUX2_X1 port map( A => SIG_in(16), B => N15, S => n2_port, Z => 
                           SIG_out(16));
   U22 : MUX2_X1 port map( A => SIG_in(17), B => N16, S => n2_port, Z => 
                           SIG_out(17));
   U23 : MUX2_X1 port map( A => SIG_in(18), B => N17, S => n2_port, Z => 
                           SIG_out(18));
   U24 : MUX2_X1 port map( A => SIG_in(19), B => N18, S => n2_port, Z => 
                           SIG_out(19));
   U25 : MUX2_X1 port map( A => SIG_in(20), B => N19, S => n2_port, Z => 
                           SIG_out(20));
   U26 : MUX2_X1 port map( A => SIG_in(21), B => N20, S => n2_port, Z => 
                           SIG_out(21));
   U27 : MUX2_X1 port map( A => SIG_in(22), B => N21, S => n2_port, Z => 
                           SIG_out(22));
   U28 : MUX2_X1 port map( A => SIG_in(23), B => N22, S => n2_port, Z => 
                           SIG_out(23));
   U29 : MUX2_X1 port map( A => SIG_in(24), B => N23, S => n2_port, Z => 
                           SIG_out(24));
   U30 : MUX2_X1 port map( A => SIG_in(25), B => N24, S => n2_port, Z => 
                           SIG_out(25));
   U31 : MUX2_X1 port map( A => SIG_in(26), B => N25, S => n2_port, Z => 
                           SIG_out(26));
   U32 : MUX2_X1 port map( A => SIG_in(27), B => N26, S => n1, Z => SIG_out(27)
                           );

end SYN_FPround;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPnormalize_SIG_width28_0 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0));

end FPnormalize_SIG_width28_0;

architecture SYN_FPnormalize of FPnormalize_SIG_width28_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17 : std_logic;

begin
   
   SIG_out(27) <= '0';
   U2 : INV_X1 port map( A => n2, ZN => n1);
   U3 : XNOR2_X1 port map( A => EXP_in(6), B => n14, ZN => EXP_out(6));
   U4 : INV_X1 port map( A => SIG_in(27), ZN => n2);
   U5 : XOR2_X1 port map( A => EXP_in(0), B => SIG_in(27), Z => EXP_out(0));
   U6 : INV_X1 port map( A => EXP_in(0), ZN => n3);
   U7 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => n4);
   U8 : XOR2_X1 port map( A => EXP_in(1), B => n4, Z => EXP_out(1));
   U9 : NAND3_X1 port map( A1 => EXP_in(1), A2 => n1, A3 => EXP_in(0), ZN => n5
                           );
   U10 : INV_X1 port map( A => n5, ZN => n8);
   U11 : XOR2_X1 port map( A => EXP_in(2), B => n8, Z => EXP_out(2));
   U12 : INV_X1 port map( A => EXP_in(2), ZN => n6);
   U13 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => n7);
   U14 : XOR2_X1 port map( A => EXP_in(3), B => n7, Z => EXP_out(3));
   U15 : NAND3_X1 port map( A1 => EXP_in(3), A2 => EXP_in(2), A3 => n8, ZN => 
                           n9);
   U16 : INV_X1 port map( A => n9, ZN => n12);
   U17 : XOR2_X1 port map( A => EXP_in(4), B => n12, Z => EXP_out(4));
   U18 : INV_X1 port map( A => EXP_in(4), ZN => n10);
   U19 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n11);
   U20 : XOR2_X1 port map( A => EXP_in(5), B => n11, Z => EXP_out(5));
   U21 : NAND3_X1 port map( A1 => EXP_in(5), A2 => EXP_in(4), A3 => n12, ZN => 
                           n14);
   U22 : INV_X1 port map( A => EXP_in(6), ZN => n13);
   U23 : NOR2_X1 port map( A1 => n14, A2 => n13, ZN => n15);
   U24 : XOR2_X1 port map( A => EXP_in(7), B => n15, Z => EXP_out(7));
   U25 : OAI21_X1 port map( B1 => SIG_in(1), B2 => n2, A => SIG_in(0), ZN => 
                           n16);
   U26 : INV_X1 port map( A => n16, ZN => SIG_out(0));
   U27 : MUX2_X1 port map( A => SIG_in(1), B => SIG_in(2), S => n1, Z => 
                           SIG_out(1));
   U28 : MUX2_X1 port map( A => SIG_in(2), B => SIG_in(3), S => n1, Z => 
                           SIG_out(2));
   U29 : MUX2_X1 port map( A => SIG_in(3), B => SIG_in(4), S => n1, Z => 
                           SIG_out(3));
   U30 : MUX2_X1 port map( A => SIG_in(4), B => SIG_in(5), S => n1, Z => 
                           SIG_out(4));
   U31 : MUX2_X1 port map( A => SIG_in(5), B => SIG_in(6), S => n1, Z => 
                           SIG_out(5));
   U32 : MUX2_X1 port map( A => SIG_in(6), B => SIG_in(7), S => n1, Z => 
                           SIG_out(6));
   U33 : MUX2_X1 port map( A => SIG_in(7), B => SIG_in(8), S => n1, Z => 
                           SIG_out(7));
   U34 : MUX2_X1 port map( A => SIG_in(8), B => SIG_in(9), S => n1, Z => 
                           SIG_out(8));
   U35 : MUX2_X1 port map( A => SIG_in(9), B => SIG_in(10), S => n1, Z => 
                           SIG_out(9));
   U36 : MUX2_X1 port map( A => SIG_in(10), B => SIG_in(11), S => n1, Z => 
                           SIG_out(10));
   U37 : MUX2_X1 port map( A => SIG_in(11), B => SIG_in(12), S => n1, Z => 
                           SIG_out(11));
   U38 : MUX2_X1 port map( A => SIG_in(12), B => SIG_in(13), S => n1, Z => 
                           SIG_out(12));
   U39 : MUX2_X1 port map( A => SIG_in(13), B => SIG_in(14), S => SIG_in(27), Z
                           => SIG_out(13));
   U40 : MUX2_X1 port map( A => SIG_in(14), B => SIG_in(15), S => SIG_in(27), Z
                           => SIG_out(14));
   U41 : MUX2_X1 port map( A => SIG_in(15), B => SIG_in(16), S => SIG_in(27), Z
                           => SIG_out(15));
   U42 : MUX2_X1 port map( A => SIG_in(16), B => SIG_in(17), S => SIG_in(27), Z
                           => SIG_out(16));
   U43 : MUX2_X1 port map( A => SIG_in(17), B => SIG_in(18), S => SIG_in(27), Z
                           => SIG_out(17));
   U44 : MUX2_X1 port map( A => SIG_in(18), B => SIG_in(19), S => SIG_in(27), Z
                           => SIG_out(18));
   U45 : MUX2_X1 port map( A => SIG_in(19), B => SIG_in(20), S => SIG_in(27), Z
                           => SIG_out(19));
   U46 : MUX2_X1 port map( A => SIG_in(20), B => SIG_in(21), S => SIG_in(27), Z
                           => SIG_out(20));
   U47 : MUX2_X1 port map( A => SIG_in(21), B => SIG_in(22), S => SIG_in(27), Z
                           => SIG_out(21));
   U48 : MUX2_X1 port map( A => SIG_in(22), B => SIG_in(23), S => SIG_in(27), Z
                           => SIG_out(22));
   U49 : MUX2_X1 port map( A => SIG_in(23), B => SIG_in(24), S => SIG_in(27), Z
                           => SIG_out(23));
   U50 : MUX2_X1 port map( A => SIG_in(24), B => SIG_in(25), S => SIG_in(27), Z
                           => SIG_out(24));
   U51 : MUX2_X1 port map( A => SIG_in(25), B => SIG_in(26), S => SIG_in(27), Z
                           => SIG_out(25));
   U52 : INV_X1 port map( A => SIG_in(26), ZN => n17);
   U53 : NAND2_X1 port map( A1 => n17, A2 => n2, ZN => SIG_out(26));

end SYN_FPnormalize;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MBE is

   port( A, B : in std_logic_vector (31 downto 0);  C : out std_logic_vector 
         (63 downto 0));

end MBE;

architecture SYN_beh of MBE is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (63 downto 0);  Cout : out std_logic);
   end component;
   
   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_1
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_2
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_3
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_4
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_5
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_6
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_7
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_8
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_9
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_10
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_11
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_12
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_345
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_346
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_347
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_348
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_349
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_350
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_351
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_352
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_353
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_354
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_355
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_356
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_357
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_358
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_359
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_360
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_361
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_362
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_363
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_364
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_365
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_378
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_13
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_14
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_15
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_381
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_382
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_383
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_384
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_385
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_386
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_388
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_389
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_390
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_16
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_17
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_18
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_421
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_422
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_423
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_424
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_425
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_426
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_427
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_428
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_19
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_20
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_21
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_465
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_466
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_467
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_468
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_469
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_470
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_471
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_472
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_473
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_474
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_475
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_476
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_477
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_478
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_479
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_480
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_482
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_22
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_23
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_24
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_485
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_486
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_487
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_488
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_489
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_490
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_491
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_492
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_493
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_25
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_26
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_27
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_512
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_513
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_514
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_515
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_516
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_517
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_518
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_519
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_520
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_521
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_522
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_523
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_524
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_525
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_526
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_527
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_528
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_529
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_530
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_531
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_532
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_533
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_534
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_535
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_536
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_28
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_29
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_30
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_537
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_538
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_539
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_540
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_541
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_542
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_543
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_544
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_545
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_546
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_547
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_548
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_549
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_550
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_551
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_552
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_553
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_554
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_555
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_556
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_557
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_558
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_559
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_560
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_561
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_562
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_563
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_564
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_565
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_566
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_567
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_568
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_31
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_32
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_33
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_569
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_570
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_571
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_572
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_34
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_35
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_36
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_573
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_574
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_575
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_576
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_577
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_578
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_579
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_580
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_37
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_38
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_39
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_581
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_582
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_583
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_584
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_585
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_586
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_587
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_588
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_589
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_590
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_591
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_592
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_40
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_41
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_42
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_593
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_594
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_595
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_596
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_597
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_598
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_599
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_600
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_601
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_602
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_603
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_604
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_605
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_606
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_607
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_43
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_0
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component ENC_1
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_2
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_3
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_4
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_5
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_6
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_7
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_8
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_9
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_10
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_11
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_12
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_13
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_14
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_15
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_16
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   component ENC_0
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, q_0_0_32_port, q_0_0_31_port, 
      q_0_0_30_port, q_0_0_29_port, q_0_0_28_port, q_0_0_27_port, q_0_0_26_port
      , q_0_0_25_port, q_0_0_24_port, q_0_0_23_port, q_0_0_22_port, 
      q_0_0_21_port, q_0_0_20_port, q_0_0_19_port, q_0_0_18_port, q_0_0_17_port
      , q_0_0_16_port, q_0_0_15_port, q_0_0_14_port, q_0_0_13_port, 
      q_0_0_12_port, q_0_0_11_port, q_0_0_10_port, q_0_0_9_port, q_0_0_8_port, 
      q_0_0_7_port, q_0_0_6_port, q_0_0_5_port, q_0_0_4_port, q_0_0_3_port, 
      q_0_0_2_port, q_0_0_1_port, q_0_0_0_port, q_0_8_50_port, q_0_8_49_port, 
      q_0_8_48_port, q_0_8_47_port, q_0_8_46_port, q_0_8_45_port, q_0_8_44_port
      , q_0_8_43_port, q_0_8_42_port, q_0_8_41_port, q_0_8_40_port, 
      q_0_8_39_port, q_0_8_38_port, q_0_8_37_port, q_0_8_36_port, q_0_8_35_port
      , q_0_8_34_port, q_0_8_33_port, q_0_8_32_port, q_0_8_31_port, 
      q_0_8_30_port, q_0_8_29_port, q_0_8_28_port, q_0_8_27_port, q_0_8_26_port
      , q_0_8_25_port, q_0_8_24_port, q_0_8_23_port, q_0_8_22_port, 
      q_0_8_21_port, q_0_8_20_port, q_0_8_19_port, q_0_8_18_port, q_0_8_17_port
      , q_0_8_16_port, q_0_7_52_port, q_0_7_51_port, q_0_7_50_port, 
      q_0_7_49_port, q_0_7_48_port, q_0_7_47_port, q_0_7_46_port, q_0_7_45_port
      , q_0_7_44_port, q_0_7_43_port, q_0_7_42_port, q_0_7_41_port, 
      q_0_7_40_port, q_0_7_39_port, q_0_7_38_port, q_0_7_37_port, q_0_7_36_port
      , q_0_7_35_port, q_0_7_34_port, q_0_7_33_port, q_0_7_32_port, 
      q_0_7_31_port, q_0_7_30_port, q_0_7_29_port, q_0_7_28_port, q_0_7_27_port
      , q_0_7_26_port, q_0_7_25_port, q_0_7_24_port, q_0_7_23_port, 
      q_0_7_22_port, q_0_7_21_port, q_0_7_20_port, q_0_7_19_port, q_0_7_18_port
      , q_0_7_17_port, q_0_7_16_port, q_0_7_15_port, q_0_7_14_port, 
      q_0_6_54_port, q_0_6_53_port, q_0_6_52_port, q_0_6_51_port, q_0_6_50_port
      , q_0_6_49_port, q_0_6_48_port, q_0_6_47_port, q_0_6_46_port, 
      q_0_6_45_port, q_0_6_44_port, q_0_6_43_port, q_0_6_42_port, q_0_6_41_port
      , q_0_6_40_port, q_0_6_39_port, q_0_6_38_port, q_0_6_37_port, 
      q_0_6_36_port, q_0_6_35_port, q_0_6_34_port, q_0_6_33_port, q_0_6_32_port
      , q_0_6_31_port, q_0_6_30_port, q_0_6_29_port, q_0_6_28_port, 
      q_0_6_27_port, q_0_6_26_port, q_0_6_25_port, q_0_6_24_port, q_0_6_23_port
      , q_0_6_22_port, q_0_6_21_port, q_0_6_20_port, q_0_6_19_port, 
      q_0_6_18_port, q_0_6_17_port, q_0_6_16_port, q_0_6_15_port, q_0_6_14_port
      , q_0_6_13_port, q_0_6_12_port, q_0_5_56_port, q_0_5_55_port, 
      q_0_5_54_port, q_0_5_53_port, q_0_5_52_port, q_0_5_51_port, q_0_5_50_port
      , q_0_5_49_port, q_0_5_48_port, q_0_5_47_port, q_0_5_46_port, 
      q_0_5_45_port, q_0_5_44_port, q_0_5_43_port, q_0_5_42_port, q_0_5_41_port
      , q_0_5_40_port, q_0_5_39_port, q_0_5_38_port, q_0_5_37_port, 
      q_0_5_36_port, q_0_5_35_port, q_0_5_34_port, q_0_5_33_port, q_0_5_32_port
      , q_0_5_31_port, q_0_5_30_port, q_0_5_29_port, q_0_5_28_port, 
      q_0_5_27_port, q_0_5_26_port, q_0_5_25_port, q_0_5_24_port, q_0_5_23_port
      , q_0_5_22_port, q_0_5_21_port, q_0_5_20_port, q_0_5_19_port, 
      q_0_5_18_port, q_0_5_17_port, q_0_5_16_port, q_0_5_15_port, q_0_5_14_port
      , q_0_5_13_port, q_0_5_12_port, q_0_5_11_port, q_0_5_10_port, 
      q_0_4_58_port, q_0_4_57_port, q_0_4_56_port, q_0_4_55_port, q_0_4_54_port
      , q_0_4_53_port, q_0_4_52_port, q_0_4_51_port, q_0_4_50_port, 
      q_0_4_49_port, q_0_4_48_port, q_0_4_47_port, q_0_4_46_port, q_0_4_45_port
      , q_0_4_44_port, q_0_4_43_port, q_0_4_42_port, q_0_4_41_port, 
      q_0_4_40_port, q_0_4_39_port, q_0_4_38_port, q_0_4_37_port, q_0_4_36_port
      , q_0_4_35_port, q_0_4_34_port, q_0_4_33_port, q_0_4_32_port, 
      q_0_4_31_port, q_0_4_30_port, q_0_4_29_port, q_0_4_28_port, q_0_4_27_port
      , q_0_4_26_port, q_0_4_25_port, q_0_4_24_port, q_0_4_23_port, 
      q_0_4_22_port, q_0_4_21_port, q_0_4_20_port, q_0_4_19_port, q_0_4_18_port
      , q_0_4_17_port, q_0_4_16_port, q_0_4_15_port, q_0_4_14_port, 
      q_0_4_13_port, q_0_4_12_port, q_0_4_11_port, q_0_4_10_port, q_0_4_9_port,
      q_0_4_8_port, q_0_3_60_port, q_0_3_59_port, q_0_3_58_port, q_0_3_57_port,
      q_0_3_56_port, q_0_3_55_port, q_0_3_54_port, q_0_3_53_port, q_0_3_52_port
      , q_0_3_51_port, q_0_3_50_port, q_0_3_49_port, q_0_3_48_port, 
      q_0_3_47_port, q_0_3_46_port, q_0_3_45_port, q_0_3_44_port, q_0_3_43_port
      , q_0_3_42_port, q_0_3_41_port, q_0_3_40_port, q_0_3_39_port, 
      q_0_3_38_port, q_0_3_37_port, q_0_3_36_port, q_0_3_35_port, q_0_3_34_port
      , q_0_3_33_port, q_0_3_32_port, q_0_3_31_port, q_0_3_30_port, 
      q_0_3_29_port, q_0_3_28_port, q_0_3_27_port, q_0_3_26_port, q_0_3_25_port
      , q_0_3_24_port, q_0_3_23_port, q_0_3_22_port, q_0_3_21_port, 
      q_0_3_20_port, q_0_3_19_port, q_0_3_18_port, q_0_3_17_port, q_0_3_16_port
      , q_0_3_15_port, q_0_3_14_port, q_0_3_13_port, q_0_3_12_port, 
      q_0_3_11_port, q_0_3_10_port, q_0_3_9_port, q_0_3_8_port, q_0_3_7_port, 
      q_0_3_6_port, q_0_2_62_port, q_0_2_61_port, q_0_2_60_port, q_0_2_59_port,
      q_0_2_58_port, q_0_2_57_port, q_0_2_56_port, q_0_2_55_port, q_0_2_54_port
      , q_0_2_53_port, q_0_2_52_port, q_0_2_51_port, q_0_2_50_port, 
      q_0_2_49_port, q_0_2_48_port, q_0_2_47_port, q_0_2_46_port, q_0_2_45_port
      , q_0_2_44_port, q_0_2_43_port, q_0_2_42_port, q_0_2_41_port, 
      q_0_2_40_port, q_0_2_39_port, q_0_2_38_port, q_0_2_37_port, q_0_2_36_port
      , q_0_2_35_port, q_0_2_34_port, q_0_2_33_port, q_0_2_32_port, 
      q_0_2_31_port, q_0_2_30_port, q_0_2_29_port, q_0_2_28_port, q_0_2_27_port
      , q_0_2_26_port, q_0_2_25_port, q_0_2_24_port, q_0_2_23_port, 
      q_0_2_22_port, q_0_2_21_port, q_0_2_20_port, q_0_2_19_port, q_0_2_18_port
      , q_0_2_17_port, q_0_2_16_port, q_0_2_15_port, q_0_2_14_port, 
      q_0_2_13_port, q_0_2_12_port, q_0_2_11_port, q_0_2_10_port, q_0_2_9_port,
      q_0_2_8_port, q_0_2_7_port, q_0_2_6_port, q_0_2_5_port, q_0_2_4_port, 
      q_0_1_63_port, q_0_1_62_port, q_0_1_61_port, q_0_1_60_port, q_0_1_59_port
      , q_0_1_58_port, q_0_1_57_port, q_0_1_56_port, q_0_1_55_port, 
      q_0_1_54_port, q_0_1_53_port, q_0_1_52_port, q_0_1_51_port, q_0_1_50_port
      , q_0_1_49_port, q_0_1_48_port, q_0_1_47_port, q_0_1_46_port, 
      q_0_1_45_port, q_0_1_44_port, q_0_1_43_port, q_0_1_42_port, q_0_1_41_port
      , q_0_1_40_port, q_0_1_39_port, q_0_1_38_port, q_0_1_37_port, 
      q_0_1_36_port, q_0_1_34_port, q_0_1_33_port, q_0_1_32_port, q_0_1_31_port
      , q_0_1_30_port, q_0_1_29_port, q_0_1_28_port, q_0_1_27_port, 
      q_0_1_26_port, q_0_1_25_port, q_0_1_24_port, q_0_1_23_port, q_0_1_22_port
      , q_0_1_21_port, q_0_1_20_port, q_0_1_19_port, q_0_1_18_port, 
      q_0_1_17_port, q_0_1_16_port, q_0_1_15_port, q_0_1_14_port, q_0_1_13_port
      , q_0_1_12_port, q_0_1_11_port, q_0_1_10_port, q_0_1_9_port, q_0_1_8_port
      , q_0_1_7_port, q_0_1_6_port, q_0_1_5_port, q_0_1_4_port, q_0_1_3_port, 
      q_0_1_2_port, q_0_16_35_port, q_0_16_34_port, q_0_16_33_port, 
      q_0_16_32_port, q_0_15_36_port, q_0_15_35_port, q_0_15_34_port, 
      q_0_15_33_port, q_0_15_32_port, q_0_15_31_port, q_0_15_30_port, 
      q_0_14_38_port, q_0_14_37_port, q_0_14_36_port, q_0_14_35_port, 
      q_0_14_34_port, q_0_14_33_port, q_0_14_32_port, q_0_14_31_port, 
      q_0_14_30_port, q_0_14_29_port, q_0_14_28_port, q_0_13_40_port, 
      q_0_13_39_port, q_0_13_38_port, q_0_13_37_port, q_0_13_36_port, 
      q_0_13_35_port, q_0_13_34_port, q_0_13_33_port, q_0_13_32_port, 
      q_0_13_31_port, q_0_13_30_port, q_0_13_29_port, q_0_13_28_port, 
      q_0_13_27_port, q_0_13_26_port, q_0_12_42_port, q_0_12_41_port, 
      q_0_12_40_port, q_0_12_39_port, q_0_12_38_port, q_0_12_37_port, 
      q_0_12_36_port, q_0_12_35_port, q_0_12_34_port, q_0_12_33_port, 
      q_0_12_32_port, q_0_12_31_port, q_0_12_30_port, q_0_12_29_port, 
      q_0_12_28_port, q_0_12_27_port, q_0_12_26_port, q_0_12_25_port, 
      q_0_12_24_port, q_0_11_44_port, q_0_11_43_port, q_0_11_42_port, 
      q_0_11_41_port, q_0_11_40_port, q_0_11_39_port, q_0_11_38_port, 
      q_0_11_37_port, q_0_11_36_port, q_0_11_35_port, q_0_11_34_port, 
      q_0_11_33_port, q_0_11_32_port, q_0_11_31_port, q_0_11_30_port, 
      q_0_11_29_port, q_0_11_28_port, q_0_11_27_port, q_0_11_26_port, 
      q_0_11_25_port, q_0_11_24_port, q_0_11_23_port, q_0_11_22_port, 
      q_0_10_46_port, q_0_10_45_port, q_0_10_44_port, q_0_10_43_port, 
      q_0_10_42_port, q_0_10_41_port, q_0_10_40_port, q_0_10_39_port, 
      q_0_10_38_port, q_0_10_37_port, q_0_10_36_port, q_0_10_35_port, 
      q_0_10_34_port, q_0_10_33_port, q_0_10_32_port, q_0_10_31_port, 
      q_0_10_30_port, q_0_10_29_port, q_0_10_28_port, q_0_10_27_port, 
      q_0_10_26_port, q_0_10_25_port, q_0_10_24_port, q_0_10_23_port, 
      q_0_10_22_port, q_0_10_21_port, q_0_10_20_port, q_0_9_48_port, 
      q_0_9_47_port, q_0_9_46_port, q_0_9_45_port, q_0_9_44_port, q_0_9_43_port
      , q_0_9_42_port, q_0_9_41_port, q_0_9_40_port, q_0_9_39_port, 
      q_0_9_38_port, q_0_9_37_port, q_0_9_36_port, q_0_9_35_port, q_0_9_34_port
      , q_0_9_33_port, q_0_9_32_port, q_0_9_31_port, q_0_9_30_port, 
      q_0_9_29_port, q_0_9_28_port, q_0_9_27_port, q_0_9_26_port, q_0_9_25_port
      , q_0_9_24_port, q_0_9_23_port, q_0_9_22_port, q_0_9_21_port, 
      q_0_9_20_port, q_0_9_19_port, q_0_9_18_port, q_1_1_42_port, q_1_1_41_port
      , q_1_1_40_port, q_1_1_39_port, q_1_1_38_port, q_1_1_37_port, 
      q_1_1_36_port, q_1_1_35_port, q_1_1_34_port, q_1_1_33_port, q_1_1_32_port
      , q_1_1_31_port, q_1_1_30_port, q_1_1_29_port, q_1_1_28_port, 
      q_1_1_27_port, q_1_1_26_port, q_1_1_25_port, q_1_0_43_port, q_1_0_42_port
      , q_1_0_41_port, q_1_0_40_port, q_1_0_39_port, q_1_0_38_port, 
      q_1_0_37_port, q_1_0_36_port, q_1_0_35_port, q_1_0_34_port, q_1_0_33_port
      , q_1_0_32_port, q_1_0_31_port, q_1_0_30_port, q_1_0_29_port, 
      q_1_0_28_port, q_1_0_27_port, q_1_0_26_port, q_1_0_25_port, q_1_0_24_port
      , q_1_7_36_port, q_1_7_35_port, q_1_7_34_port, q_1_7_33_port, 
      q_1_7_32_port, q_1_7_31_port, q_1_6_37_port, q_1_6_36_port, q_1_6_35_port
      , q_1_6_34_port, q_1_6_33_port, q_1_6_32_port, q_1_6_31_port, 
      q_1_6_30_port, q_1_5_38_port, q_1_5_37_port, q_1_5_36_port, q_1_5_35_port
      , q_1_5_34_port, q_1_5_33_port, q_1_5_32_port, q_1_5_31_port, 
      q_1_5_30_port, q_1_5_29_port, q_1_4_39_port, q_1_4_38_port, q_1_4_37_port
      , q_1_4_36_port, q_1_4_35_port, q_1_4_34_port, q_1_4_33_port, 
      q_1_4_32_port, q_1_4_31_port, q_1_4_30_port, q_1_4_29_port, q_1_4_28_port
      , q_1_3_40_port, q_1_3_39_port, q_1_3_38_port, q_1_3_37_port, 
      q_1_3_36_port, q_1_3_35_port, q_1_3_34_port, q_1_3_33_port, q_1_3_32_port
      , q_1_3_31_port, q_1_3_30_port, q_1_3_29_port, q_1_3_28_port, 
      q_1_3_27_port, q_1_2_41_port, q_1_2_40_port, q_1_2_39_port, q_1_2_38_port
      , q_1_2_37_port, q_1_2_36_port, q_1_2_35_port, q_1_2_34_port, 
      q_1_2_33_port, q_1_2_32_port, q_1_2_31_port, q_1_2_30_port, q_1_2_29_port
      , q_1_2_28_port, q_1_2_27_port, q_1_2_26_port, q_2_2_49_port, 
      q_2_2_48_port, q_2_2_47_port, q_2_2_46_port, q_2_2_45_port, q_2_2_44_port
      , q_2_2_43_port, q_2_2_42_port, q_2_2_41_port, q_2_2_40_port, 
      q_2_2_39_port, q_2_2_38_port, q_2_2_37_port, q_2_2_36_port, q_2_2_35_port
      , q_2_2_34_port, q_2_2_33_port, q_2_2_32_port, q_2_2_31_port, 
      q_2_2_30_port, q_2_2_29_port, q_2_2_28_port, q_2_2_27_port, q_2_2_26_port
      , q_2_2_25_port, q_2_2_24_port, q_2_2_23_port, q_2_2_22_port, 
      q_2_2_21_port, q_2_2_20_port, q_2_2_19_port, q_2_2_18_port, q_2_1_50_port
      , q_2_1_49_port, q_2_1_48_port, q_2_1_47_port, q_2_1_46_port, 
      q_2_1_45_port, q_2_1_44_port, q_2_1_43_port, q_2_1_42_port, q_2_1_41_port
      , q_2_1_40_port, q_2_1_39_port, q_2_1_38_port, q_2_1_37_port, 
      q_2_1_36_port, q_2_1_35_port, q_2_1_34_port, q_2_1_33_port, q_2_1_32_port
      , q_2_1_31_port, q_2_1_30_port, q_2_1_29_port, q_2_1_28_port, 
      q_2_1_27_port, q_2_1_26_port, q_2_1_25_port, q_2_1_24_port, q_2_1_23_port
      , q_2_1_22_port, q_2_1_21_port, q_2_1_20_port, q_2_1_19_port, 
      q_2_1_18_port, q_2_1_17_port, q_2_0_51_port, q_2_0_50_port, q_2_0_49_port
      , q_2_0_48_port, q_2_0_47_port, q_2_0_46_port, q_2_0_45_port, 
      q_2_0_44_port, q_2_0_43_port, q_2_0_42_port, q_2_0_41_port, q_2_0_40_port
      , q_2_0_39_port, q_2_0_38_port, q_2_0_37_port, q_2_0_36_port, 
      q_2_0_35_port, q_2_0_34_port, q_2_0_33_port, q_2_0_32_port, q_2_0_31_port
      , q_2_0_30_port, q_2_0_29_port, q_2_0_28_port, q_2_0_27_port, 
      q_2_0_26_port, q_2_0_25_port, q_2_0_24_port, q_2_0_23_port, q_2_0_22_port
      , q_2_0_21_port, q_2_0_20_port, q_2_0_19_port, q_2_0_18_port, 
      q_2_0_17_port, q_2_0_16_port, q_2_7_44_port, q_2_7_43_port, q_2_7_42_port
      , q_2_7_41_port, q_2_7_40_port, q_2_7_39_port, q_2_7_38_port, 
      q_2_7_37_port, q_2_7_36_port, q_2_7_35_port, q_2_7_34_port, q_2_7_33_port
      , q_2_7_32_port, q_2_7_31_port, q_2_7_30_port, q_2_7_29_port, 
      q_2_7_28_port, q_2_7_27_port, q_2_7_26_port, q_2_7_25_port, q_2_7_24_port
      , q_2_7_23_port, q_2_6_45_port, q_2_6_44_port, q_2_6_43_port, 
      q_2_6_42_port, q_2_6_41_port, q_2_6_40_port, q_2_6_39_port, q_2_6_38_port
      , q_2_6_37_port, q_2_6_36_port, q_2_6_35_port, q_2_6_34_port, 
      q_2_6_33_port, q_2_6_32_port, q_2_6_31_port, q_2_6_30_port, q_2_6_29_port
      , q_2_6_28_port, q_2_6_27_port, q_2_6_26_port, q_2_6_25_port, 
      q_2_6_24_port, q_2_6_23_port, q_2_6_22_port, q_2_5_46_port, q_2_5_45_port
      , q_2_5_44_port, q_2_5_43_port, q_2_5_42_port, q_2_5_41_port, 
      q_2_5_40_port, q_2_5_39_port, q_2_5_38_port, q_2_5_37_port, q_2_5_36_port
      , q_2_5_35_port, q_2_5_34_port, q_2_5_33_port, q_2_5_32_port, 
      q_2_5_31_port, q_2_5_30_port, q_2_5_29_port, q_2_5_28_port, q_2_5_27_port
      , q_2_5_26_port, q_2_5_25_port, q_2_5_24_port, q_2_5_23_port, 
      q_2_5_22_port, q_2_5_21_port, q_2_4_47_port, q_2_4_46_port, q_2_4_45_port
      , q_2_4_44_port, q_2_4_43_port, q_2_4_42_port, q_2_4_41_port, 
      q_2_4_40_port, q_2_4_39_port, q_2_4_38_port, q_2_4_37_port, q_2_4_36_port
      , q_2_4_35_port, q_2_4_34_port, q_2_4_33_port, q_2_4_32_port, 
      q_2_4_31_port, q_2_4_30_port, q_2_4_29_port, q_2_4_28_port, q_2_4_27_port
      , q_2_4_26_port, q_2_4_25_port, q_2_4_24_port, q_2_4_23_port, 
      q_2_4_22_port, q_2_4_21_port, q_2_4_20_port, q_2_3_48_port, q_2_3_47_port
      , q_2_3_46_port, q_2_3_45_port, q_2_3_44_port, q_2_3_43_port, 
      q_2_3_42_port, q_2_3_41_port, q_2_3_40_port, q_2_3_39_port, q_2_3_38_port
      , q_2_3_37_port, q_2_3_36_port, q_2_3_35_port, q_2_3_34_port, 
      q_2_3_33_port, q_2_3_32_port, q_2_3_31_port, q_2_3_30_port, q_2_3_29_port
      , q_2_3_28_port, q_2_3_27_port, q_2_3_26_port, q_2_3_25_port, 
      q_2_3_24_port, q_2_3_23_port, q_2_3_22_port, q_2_3_21_port, q_2_3_20_port
      , q_2_3_19_port, q_3_3_54_port, q_3_3_53_port, q_3_3_52_port, 
      q_3_3_51_port, q_3_3_50_port, q_3_3_49_port, q_3_3_48_port, q_3_3_47_port
      , q_3_3_46_port, q_3_3_45_port, q_3_3_44_port, q_3_3_43_port, 
      q_3_3_42_port, q_3_3_41_port, q_3_3_40_port, q_3_3_39_port, q_3_3_38_port
      , q_3_3_37_port, q_3_3_36_port, q_3_3_35_port, q_3_3_34_port, 
      q_3_3_33_port, q_3_3_32_port, q_3_3_31_port, q_3_3_30_port, q_3_3_29_port
      , q_3_3_28_port, q_3_3_27_port, q_3_3_26_port, q_3_3_25_port, 
      q_3_3_24_port, q_3_3_23_port, q_3_3_22_port, q_3_3_21_port, q_3_3_20_port
      , q_3_3_19_port, q_3_3_18_port, q_3_3_17_port, q_3_3_16_port, 
      q_3_3_15_port, q_3_3_14_port, q_3_3_13_port, q_3_2_55_port, q_3_2_54_port
      , q_3_2_53_port, q_3_2_52_port, q_3_2_51_port, q_3_2_50_port, 
      q_3_2_49_port, q_3_2_48_port, q_3_2_47_port, q_3_2_46_port, q_3_2_45_port
      , q_3_2_44_port, q_3_2_43_port, q_3_2_42_port, q_3_2_41_port, 
      q_3_2_40_port, q_3_2_39_port, q_3_2_38_port, q_3_2_37_port, q_3_2_36_port
      , q_3_2_35_port, q_3_2_34_port, q_3_2_33_port, q_3_2_32_port, 
      q_3_2_31_port, q_3_2_30_port, q_3_2_29_port, q_3_2_28_port, q_3_2_27_port
      , q_3_2_26_port, q_3_2_25_port, q_3_2_24_port, q_3_2_23_port, 
      q_3_2_22_port, q_3_2_21_port, q_3_2_20_port, q_3_2_19_port, q_3_2_18_port
      , q_3_2_17_port, q_3_2_16_port, q_3_2_15_port, q_3_2_14_port, 
      q_3_2_13_port, q_3_2_12_port, q_3_1_56_port, q_3_1_55_port, q_3_1_54_port
      , q_3_1_53_port, q_3_1_52_port, q_3_1_51_port, q_3_1_50_port, 
      q_3_1_49_port, q_3_1_48_port, q_3_1_47_port, q_3_1_46_port, q_3_1_45_port
      , q_3_1_44_port, q_3_1_43_port, q_3_1_42_port, q_3_1_41_port, 
      q_3_1_40_port, q_3_1_39_port, q_3_1_38_port, q_3_1_37_port, q_3_1_36_port
      , q_3_1_35_port, q_3_1_34_port, q_3_1_33_port, q_3_1_32_port, 
      q_3_1_31_port, q_3_1_30_port, q_3_1_29_port, q_3_1_28_port, q_3_1_27_port
      , q_3_1_26_port, q_3_1_25_port, q_3_1_24_port, q_3_1_23_port, 
      q_3_1_22_port, q_3_1_21_port, q_3_1_20_port, q_3_1_19_port, q_3_1_18_port
      , q_3_1_17_port, q_3_1_16_port, q_3_1_15_port, q_3_1_14_port, 
      q_3_1_13_port, q_3_1_12_port, q_3_1_11_port, q_3_0_57_port, q_3_0_56_port
      , q_3_0_55_port, q_3_0_54_port, q_3_0_53_port, q_3_0_52_port, 
      q_3_0_51_port, q_3_0_50_port, q_3_0_49_port, q_3_0_48_port, q_3_0_47_port
      , q_3_0_46_port, q_3_0_45_port, q_3_0_44_port, q_3_0_43_port, 
      q_3_0_42_port, q_3_0_41_port, q_3_0_40_port, q_3_0_39_port, q_3_0_38_port
      , q_3_0_37_port, q_3_0_36_port, q_3_0_35_port, q_3_0_34_port, 
      q_3_0_33_port, q_3_0_32_port, q_3_0_31_port, q_3_0_30_port, q_3_0_29_port
      , q_3_0_28_port, q_3_0_27_port, q_3_0_26_port, q_3_0_25_port, 
      q_3_0_24_port, q_3_0_23_port, q_3_0_22_port, q_3_0_21_port, q_3_0_20_port
      , q_3_0_19_port, q_3_0_18_port, q_3_0_17_port, q_3_0_16_port, 
      q_3_0_15_port, q_3_0_14_port, q_3_0_13_port, q_3_0_12_port, q_3_0_11_port
      , q_3_0_10_port, q_3_5_52_port, q_3_5_51_port, q_3_5_50_port, 
      q_3_5_49_port, q_3_5_48_port, q_3_5_47_port, q_3_5_46_port, q_3_5_45_port
      , q_3_5_44_port, q_3_5_43_port, q_3_5_42_port, q_3_5_41_port, 
      q_3_5_40_port, q_3_5_39_port, q_3_5_38_port, q_3_5_37_port, q_3_5_36_port
      , q_3_5_35_port, q_3_5_34_port, q_3_5_33_port, q_3_5_32_port, 
      q_3_5_31_port, q_3_5_30_port, q_3_5_29_port, q_3_5_28_port, q_3_5_27_port
      , q_3_5_26_port, q_3_5_25_port, q_3_5_24_port, q_3_5_23_port, 
      q_3_5_22_port, q_3_5_21_port, q_3_5_20_port, q_3_5_19_port, q_3_5_18_port
      , q_3_5_17_port, q_3_5_16_port, q_3_5_15_port, q_3_4_53_port, 
      q_3_4_52_port, q_3_4_51_port, q_3_4_50_port, q_3_4_49_port, q_3_4_48_port
      , q_3_4_47_port, q_3_4_46_port, q_3_4_45_port, q_3_4_44_port, 
      q_3_4_43_port, q_3_4_42_port, q_3_4_41_port, q_3_4_40_port, q_3_4_39_port
      , q_3_4_38_port, q_3_4_37_port, q_3_4_36_port, q_3_4_35_port, 
      q_3_4_34_port, q_3_4_33_port, q_3_4_32_port, q_3_4_31_port, q_3_4_30_port
      , q_3_4_29_port, q_3_4_28_port, q_3_4_27_port, q_3_4_26_port, 
      q_3_4_25_port, q_3_4_24_port, q_3_4_23_port, q_3_4_22_port, q_3_4_21_port
      , q_3_4_20_port, q_3_4_19_port, q_3_4_18_port, q_3_4_17_port, 
      q_3_4_16_port, q_3_4_15_port, q_3_4_14_port, q_4_2_59_port, q_4_2_58_port
      , q_4_2_57_port, q_4_2_56_port, q_4_2_55_port, q_4_2_54_port, 
      q_4_2_53_port, q_4_2_52_port, q_4_2_51_port, q_4_2_50_port, q_4_2_49_port
      , q_4_2_48_port, q_4_2_47_port, q_4_2_46_port, q_4_2_45_port, 
      q_4_2_44_port, q_4_2_43_port, q_4_2_42_port, q_4_2_41_port, q_4_2_40_port
      , q_4_2_39_port, q_4_2_38_port, q_4_2_37_port, q_4_2_36_port, 
      q_4_2_35_port, q_4_2_34_port, q_4_2_33_port, q_4_2_32_port, q_4_2_31_port
      , q_4_2_30_port, q_4_2_29_port, q_4_2_28_port, q_4_2_27_port, 
      q_4_2_26_port, q_4_2_25_port, q_4_2_24_port, q_4_2_23_port, q_4_2_22_port
      , q_4_2_21_port, q_4_2_20_port, q_4_2_19_port, q_4_2_18_port, 
      q_4_2_17_port, q_4_2_16_port, q_4_2_15_port, q_4_2_14_port, q_4_2_13_port
      , q_4_2_12_port, q_4_2_11_port, q_4_2_10_port, q_4_2_9_port, q_4_2_8_port
      , q_4_1_60_port, q_4_1_59_port, q_4_1_58_port, q_4_1_57_port, 
      q_4_1_56_port, q_4_1_55_port, q_4_1_54_port, q_4_1_53_port, q_4_1_52_port
      , q_4_1_51_port, q_4_1_50_port, q_4_1_49_port, q_4_1_48_port, 
      q_4_1_47_port, q_4_1_46_port, q_4_1_45_port, q_4_1_44_port, q_4_1_43_port
      , q_4_1_42_port, q_4_1_41_port, q_4_1_40_port, q_4_1_39_port, 
      q_4_1_38_port, q_4_1_37_port, q_4_1_36_port, q_4_1_35_port, q_4_1_34_port
      , q_4_1_33_port, q_4_1_32_port, q_4_1_31_port, q_4_1_30_port, 
      q_4_1_29_port, q_4_1_28_port, q_4_1_27_port, q_4_1_26_port, q_4_1_25_port
      , q_4_1_24_port, q_4_1_23_port, q_4_1_22_port, q_4_1_21_port, 
      q_4_1_20_port, q_4_1_19_port, q_4_1_18_port, q_4_1_17_port, q_4_1_16_port
      , q_4_1_15_port, q_4_1_14_port, q_4_1_13_port, q_4_1_12_port, 
      q_4_1_11_port, q_4_1_10_port, q_4_1_9_port, q_4_1_8_port, q_4_1_7_port, 
      q_4_0_61_port, q_4_0_60_port, q_4_0_59_port, q_4_0_58_port, q_4_0_57_port
      , q_4_0_56_port, q_4_0_55_port, q_4_0_54_port, q_4_0_53_port, 
      q_4_0_52_port, q_4_0_51_port, q_4_0_50_port, q_4_0_49_port, q_4_0_48_port
      , q_4_0_47_port, q_4_0_46_port, q_4_0_45_port, q_4_0_44_port, 
      q_4_0_43_port, q_4_0_42_port, q_4_0_41_port, q_4_0_40_port, q_4_0_39_port
      , q_4_0_38_port, q_4_0_37_port, q_4_0_36_port, q_4_0_35_port, 
      q_4_0_34_port, q_4_0_33_port, q_4_0_32_port, q_4_0_31_port, q_4_0_30_port
      , q_4_0_29_port, q_4_0_28_port, q_4_0_27_port, q_4_0_26_port, 
      q_4_0_25_port, q_4_0_24_port, q_4_0_23_port, q_4_0_22_port, q_4_0_21_port
      , q_4_0_20_port, q_4_0_19_port, q_4_0_18_port, q_4_0_17_port, 
      q_4_0_16_port, q_4_0_15_port, q_4_0_14_port, q_4_0_13_port, q_4_0_12_port
      , q_4_0_11_port, q_4_0_10_port, q_4_0_9_port, q_4_0_8_port, q_4_0_7_port,
      q_4_0_6_port, q_5_2_58_port, q_5_2_57_port, q_5_2_56_port, q_5_2_55_port,
      q_5_2_54_port, q_5_2_53_port, q_5_2_52_port, q_5_2_51_port, q_5_2_50_port
      , q_5_2_49_port, q_5_2_48_port, q_5_2_47_port, q_5_2_46_port, 
      q_5_2_45_port, q_5_2_44_port, q_5_2_43_port, q_5_2_42_port, q_5_2_41_port
      , q_5_2_40_port, q_5_2_39_port, q_5_2_38_port, q_5_2_37_port, 
      q_5_2_36_port, q_5_2_35_port, q_5_2_34_port, q_5_2_33_port, q_5_2_32_port
      , q_5_2_31_port, q_5_2_30_port, q_5_2_29_port, q_5_2_28_port, 
      q_5_2_27_port, q_5_2_26_port, q_5_2_25_port, q_5_2_24_port, q_5_2_23_port
      , q_5_2_22_port, q_5_2_21_port, q_5_2_20_port, q_5_2_19_port, 
      q_5_2_18_port, q_5_2_17_port, q_5_2_16_port, q_5_2_15_port, q_5_2_14_port
      , q_5_2_13_port, q_5_2_12_port, q_5_2_11_port, q_5_2_10_port, 
      q_5_2_9_port, q_5_1_62_port, q_5_1_61_port, q_5_1_60_port, q_5_1_59_port,
      q_5_1_58_port, q_5_1_57_port, q_5_1_56_port, q_5_1_55_port, q_5_1_54_port
      , q_5_1_53_port, q_5_1_52_port, q_5_1_51_port, q_5_1_50_port, 
      q_5_1_49_port, q_5_1_48_port, q_5_1_47_port, q_5_1_46_port, q_5_1_45_port
      , q_5_1_44_port, q_5_1_43_port, q_5_1_42_port, q_5_1_41_port, 
      q_5_1_40_port, q_5_1_39_port, q_5_1_38_port, q_5_1_37_port, q_5_1_36_port
      , q_5_1_35_port, q_5_1_34_port, q_5_1_33_port, q_5_1_32_port, 
      q_5_1_31_port, q_5_1_30_port, q_5_1_29_port, q_5_1_28_port, q_5_1_27_port
      , q_5_1_26_port, q_5_1_25_port, q_5_1_24_port, q_5_1_23_port, 
      q_5_1_22_port, q_5_1_21_port, q_5_1_20_port, q_5_1_19_port, q_5_1_18_port
      , q_5_1_17_port, q_5_1_16_port, q_5_1_15_port, q_5_1_14_port, 
      q_5_1_13_port, q_5_1_12_port, q_5_1_11_port, q_5_1_10_port, q_5_1_9_port,
      q_5_1_8_port, q_5_1_7_port, q_5_1_6_port, q_5_1_5_port, q_5_0_63_port, 
      q_5_0_62_port, q_5_0_61_port, q_5_0_60_port, q_5_0_59_port, q_5_0_58_port
      , q_5_0_57_port, q_5_0_56_port, q_5_0_55_port, q_5_0_54_port, 
      q_5_0_53_port, q_5_0_52_port, q_5_0_51_port, q_5_0_50_port, q_5_0_49_port
      , q_5_0_48_port, q_5_0_47_port, q_5_0_46_port, q_5_0_45_port, 
      q_5_0_44_port, q_5_0_43_port, q_5_0_42_port, q_5_0_41_port, q_5_0_40_port
      , q_5_0_39_port, q_5_0_38_port, q_5_0_37_port, q_5_0_36_port, 
      q_5_0_35_port, q_5_0_34_port, q_5_0_33_port, q_5_0_32_port, q_5_0_31_port
      , q_5_0_30_port, q_5_0_29_port, q_5_0_28_port, q_5_0_27_port, 
      q_5_0_26_port, q_5_0_25_port, q_5_0_24_port, q_5_0_23_port, q_5_0_22_port
      , q_5_0_21_port, q_5_0_20_port, q_5_0_19_port, q_5_0_18_port, 
      q_5_0_17_port, q_5_0_16_port, q_5_0_15_port, q_5_0_14_port, q_5_0_13_port
      , q_5_0_12_port, q_5_0_11_port, q_5_0_10_port, q_5_0_9_port, q_5_0_8_port
      , q_5_0_7_port, q_5_0_6_port, q_5_0_5_port, q_5_0_4_port, q_6_1_63_port, 
      q_6_1_62_port, q_6_1_61_port, q_6_1_60_port, q_6_1_59_port, q_6_1_58_port
      , q_6_1_57_port, q_6_1_56_port, q_6_1_55_port, q_6_1_54_port, 
      q_6_1_53_port, q_6_1_52_port, q_6_1_51_port, q_6_1_50_port, q_6_1_49_port
      , q_6_1_48_port, q_6_1_47_port, q_6_1_46_port, q_6_1_45_port, 
      q_6_1_44_port, q_6_1_43_port, q_6_1_42_port, q_6_1_41_port, q_6_1_40_port
      , q_6_1_39_port, q_6_1_38_port, q_6_1_37_port, q_6_1_36_port, 
      q_6_1_35_port, q_6_1_34_port, q_6_1_33_port, q_6_1_32_port, q_6_1_31_port
      , q_6_1_30_port, q_6_1_29_port, q_6_1_28_port, q_6_1_27_port, 
      q_6_1_26_port, q_6_1_25_port, q_6_1_24_port, q_6_1_23_port, q_6_1_22_port
      , q_6_1_21_port, q_6_1_20_port, q_6_1_19_port, q_6_1_18_port, 
      q_6_1_17_port, q_6_1_16_port, q_6_1_15_port, q_6_1_14_port, q_6_1_13_port
      , q_6_1_12_port, q_6_1_11_port, q_6_1_10_port, q_6_1_9_port, q_6_1_8_port
      , q_6_1_7_port, q_6_1_6_port, q_6_1_5_port, q_6_1_4_port, q_6_1_3_port, 
      q_6_0_63_port, q_6_0_62_port, q_6_0_61_port, q_6_0_60_port, q_6_0_59_port
      , q_6_0_58_port, q_6_0_57_port, q_6_0_56_port, q_6_0_55_port, 
      q_6_0_54_port, q_6_0_53_port, q_6_0_52_port, q_6_0_51_port, q_6_0_50_port
      , q_6_0_49_port, q_6_0_48_port, q_6_0_47_port, q_6_0_46_port, 
      q_6_0_45_port, q_6_0_44_port, q_6_0_43_port, q_6_0_42_port, q_6_0_41_port
      , q_6_0_40_port, q_6_0_39_port, q_6_0_38_port, q_6_0_37_port, 
      q_6_0_36_port, q_6_0_35_port, q_6_0_34_port, q_6_0_33_port, q_6_0_32_port
      , q_6_0_31_port, q_6_0_30_port, q_6_0_29_port, q_6_0_28_port, 
      q_6_0_27_port, q_6_0_26_port, q_6_0_25_port, q_6_0_24_port, q_6_0_23_port
      , q_6_0_22_port, q_6_0_21_port, q_6_0_20_port, q_6_0_19_port, 
      q_6_0_18_port, q_6_0_17_port, q_6_0_16_port, q_6_0_15_port, q_6_0_14_port
      , q_6_0_13_port, q_6_0_12_port, q_6_0_11_port, q_6_0_10_port, 
      q_6_0_9_port, q_6_0_8_port, q_6_0_7_port, q_6_0_6_port, q_6_0_5_port, 
      q_6_0_4_port, q_6_0_3_port, q_6_0_2_port, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n_1042, n_1043, n_1044 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   encI_1 : ENC_0 port map( b(2) => B(1), b(1) => B(0), b(0) => X_Logic0_port, 
                           A(31) => n79, A(30) => n77, A(29) => n75, A(28) => 
                           n73, A(27) => n71, A(26) => n69, A(25) => n67, A(24)
                           => n65, A(23) => n63, A(22) => n61, A(21) => n59, 
                           A(20) => n57, A(19) => n55, A(18) => n53, A(17) => 
                           n51, A(16) => n49, A(15) => n47, A(14) => n46, A(13)
                           => n44, A(12) => n42, A(11) => n40, A(10) => n38, 
                           A(9) => n36, A(8) => n34, A(7) => n32, A(6) => n30, 
                           A(5) => n28, A(4) => n26, A(3) => n24, A(2) => n22, 
                           A(1) => n20, A(0) => n18, p(32) => q_0_0_32_port, 
                           p(31) => q_0_0_31_port, p(30) => q_0_0_30_port, 
                           p(29) => q_0_0_29_port, p(28) => q_0_0_28_port, 
                           p(27) => q_0_0_27_port, p(26) => q_0_0_26_port, 
                           p(25) => q_0_0_25_port, p(24) => q_0_0_24_port, 
                           p(23) => q_0_0_23_port, p(22) => q_0_0_22_port, 
                           p(21) => q_0_0_21_port, p(20) => q_0_0_20_port, 
                           p(19) => q_0_0_19_port, p(18) => q_0_0_18_port, 
                           p(17) => q_0_0_17_port, p(16) => q_0_0_16_port, 
                           p(15) => q_0_0_15_port, p(14) => q_0_0_14_port, 
                           p(13) => q_0_0_13_port, p(12) => q_0_0_12_port, 
                           p(11) => q_0_0_11_port, p(10) => q_0_0_10_port, p(9)
                           => q_0_0_9_port, p(8) => q_0_0_8_port, p(7) => 
                           q_0_0_7_port, p(6) => q_0_0_6_port, p(5) => 
                           q_0_0_5_port, p(4) => q_0_0_4_port, p(3) => 
                           q_0_0_3_port, p(2) => q_0_0_2_port, p(1) => 
                           q_0_0_1_port, p(0) => q_0_0_0_port);
   encI_2 : ENC_16 port map( b(2) => B(3), b(1) => B(2), b(0) => B(1), A(31) =>
                           n79, A(30) => n77, A(29) => n75, A(28) => n73, A(27)
                           => n71, A(26) => n69, A(25) => n67, A(24) => n65, 
                           A(23) => n63, A(22) => n61, A(21) => n59, A(20) => 
                           n57, A(19) => n55, A(18) => n53, A(17) => n51, A(16)
                           => n49, A(15) => n47, A(14) => n45, A(13) => n43, 
                           A(12) => n41, A(11) => n39, A(10) => n37, A(9) => 
                           n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) => 
                           n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) => 
                           n19, A(0) => n17, p(32) => q_0_1_34_port, p(31) => 
                           q_0_1_33_port, p(30) => q_0_1_32_port, p(29) => 
                           q_0_1_31_port, p(28) => q_0_1_30_port, p(27) => 
                           q_0_1_29_port, p(26) => q_0_1_28_port, p(25) => 
                           q_0_1_27_port, p(24) => q_0_1_26_port, p(23) => 
                           q_0_1_25_port, p(22) => q_0_1_24_port, p(21) => 
                           q_0_1_23_port, p(20) => q_0_1_22_port, p(19) => 
                           q_0_1_21_port, p(18) => q_0_1_20_port, p(17) => 
                           q_0_1_19_port, p(16) => q_0_1_18_port, p(15) => 
                           q_0_1_17_port, p(14) => q_0_1_16_port, p(13) => 
                           q_0_1_15_port, p(12) => q_0_1_14_port, p(11) => 
                           q_0_1_13_port, p(10) => q_0_1_12_port, p(9) => 
                           q_0_1_11_port, p(8) => q_0_1_10_port, p(7) => 
                           q_0_1_9_port, p(6) => q_0_1_8_port, p(5) => 
                           q_0_1_7_port, p(4) => q_0_1_6_port, p(3) => 
                           q_0_1_5_port, p(2) => q_0_1_4_port, p(1) => 
                           q_0_1_3_port, p(0) => q_0_1_2_port);
   encI_3 : ENC_15 port map( b(2) => B(5), b(1) => B(4), b(0) => B(3), A(31) =>
                           n79, A(30) => n77, A(29) => n75, A(28) => n73, A(27)
                           => n71, A(26) => n69, A(25) => n67, A(24) => n65, 
                           A(23) => n63, A(22) => n62, A(21) => n60, A(20) => 
                           n58, A(19) => n56, A(18) => n54, A(17) => n52, A(16)
                           => n50, A(15) => n48, A(14) => n45, A(13) => n43, 
                           A(12) => n41, A(11) => n39, A(10) => n37, A(9) => 
                           n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) => 
                           n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) => 
                           n19, A(0) => n17, p(32) => q_0_1_36_port, p(31) => 
                           q_0_2_35_port, p(30) => q_0_2_34_port, p(29) => 
                           q_0_2_33_port, p(28) => q_0_2_32_port, p(27) => 
                           q_0_2_31_port, p(26) => q_0_2_30_port, p(25) => 
                           q_0_2_29_port, p(24) => q_0_2_28_port, p(23) => 
                           q_0_2_27_port, p(22) => q_0_2_26_port, p(21) => 
                           q_0_2_25_port, p(20) => q_0_2_24_port, p(19) => 
                           q_0_2_23_port, p(18) => q_0_2_22_port, p(17) => 
                           q_0_2_21_port, p(16) => q_0_2_20_port, p(15) => 
                           q_0_2_19_port, p(14) => q_0_2_18_port, p(13) => 
                           q_0_2_17_port, p(12) => q_0_2_16_port, p(11) => 
                           q_0_2_15_port, p(10) => q_0_2_14_port, p(9) => 
                           q_0_2_13_port, p(8) => q_0_2_12_port, p(7) => 
                           q_0_2_11_port, p(6) => q_0_2_10_port, p(5) => 
                           q_0_2_9_port, p(4) => q_0_2_8_port, p(3) => 
                           q_0_2_7_port, p(2) => q_0_2_6_port, p(1) => 
                           q_0_2_5_port, p(0) => q_0_2_4_port);
   encI_4 : ENC_14 port map( b(2) => B(7), b(1) => B(6), b(0) => B(5), A(31) =>
                           n79, A(30) => n77, A(29) => n75, A(28) => n73, A(27)
                           => n71, A(26) => n69, A(25) => n67, A(24) => n65, 
                           A(23) => n63, A(22) => n61, A(21) => n60, A(20) => 
                           n58, A(19) => n56, A(18) => n54, A(17) => n52, A(16)
                           => n50, A(15) => n48, A(14) => n45, A(13) => n43, 
                           A(12) => n41, A(11) => n39, A(10) => n37, A(9) => 
                           n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) => 
                           n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) => 
                           n19, A(0) => n17, p(32) => q_0_1_38_port, p(31) => 
                           q_0_1_37_port, p(30) => q_0_2_36_port, p(29) => 
                           q_0_3_35_port, p(28) => q_0_3_34_port, p(27) => 
                           q_0_3_33_port, p(26) => q_0_3_32_port, p(25) => 
                           q_0_3_31_port, p(24) => q_0_3_30_port, p(23) => 
                           q_0_3_29_port, p(22) => q_0_3_28_port, p(21) => 
                           q_0_3_27_port, p(20) => q_0_3_26_port, p(19) => 
                           q_0_3_25_port, p(18) => q_0_3_24_port, p(17) => 
                           q_0_3_23_port, p(16) => q_0_3_22_port, p(15) => 
                           q_0_3_21_port, p(14) => q_0_3_20_port, p(13) => 
                           q_0_3_19_port, p(12) => q_0_3_18_port, p(11) => 
                           q_0_3_17_port, p(10) => q_0_3_16_port, p(9) => 
                           q_0_3_15_port, p(8) => q_0_3_14_port, p(7) => 
                           q_0_3_13_port, p(6) => q_0_3_12_port, p(5) => 
                           q_0_3_11_port, p(4) => q_0_3_10_port, p(3) => 
                           q_0_3_9_port, p(2) => q_0_3_8_port, p(1) => 
                           q_0_3_7_port, p(0) => q_0_3_6_port);
   encI_5 : ENC_13 port map( b(2) => B(9), b(1) => B(8), b(0) => B(7), A(31) =>
                           n79, A(30) => n77, A(29) => n75, A(28) => n73, A(27)
                           => n71, A(26) => n69, A(25) => n67, A(24) => n65, 
                           A(23) => n63, A(22) => n61, A(21) => n60, A(20) => 
                           n57, A(19) => n55, A(18) => n54, A(17) => n52, A(16)
                           => n50, A(15) => n48, A(14) => n45, A(13) => n43, 
                           A(12) => n41, A(11) => n39, A(10) => n37, A(9) => 
                           n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) => 
                           n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) => 
                           n19, A(0) => n17, p(32) => q_0_1_40_port, p(31) => 
                           q_0_1_39_port, p(30) => q_0_2_38_port, p(29) => 
                           q_0_2_37_port, p(28) => q_0_3_36_port, p(27) => 
                           q_0_4_35_port, p(26) => q_0_4_34_port, p(25) => 
                           q_0_4_33_port, p(24) => q_0_4_32_port, p(23) => 
                           q_0_4_31_port, p(22) => q_0_4_30_port, p(21) => 
                           q_0_4_29_port, p(20) => q_0_4_28_port, p(19) => 
                           q_0_4_27_port, p(18) => q_0_4_26_port, p(17) => 
                           q_0_4_25_port, p(16) => q_0_4_24_port, p(15) => 
                           q_0_4_23_port, p(14) => q_0_4_22_port, p(13) => 
                           q_0_4_21_port, p(12) => q_0_4_20_port, p(11) => 
                           q_0_4_19_port, p(10) => q_0_4_18_port, p(9) => 
                           q_0_4_17_port, p(8) => q_0_4_16_port, p(7) => 
                           q_0_4_15_port, p(6) => q_0_4_14_port, p(5) => 
                           q_0_4_13_port, p(4) => q_0_4_12_port, p(3) => 
                           q_0_4_11_port, p(2) => q_0_4_10_port, p(1) => 
                           q_0_4_9_port, p(0) => q_0_4_8_port);
   encI_6 : ENC_12 port map( b(2) => B(11), b(1) => B(10), b(0) => B(9), A(31) 
                           => n79, A(30) => n77, A(29) => n75, A(28) => n73, 
                           A(27) => n71, A(26) => n69, A(25) => n67, A(24) => 
                           n65, A(23) => n63, A(22) => n61, A(21) => n60, A(20)
                           => n57, A(19) => n55, A(18) => n53, A(17) => n51, 
                           A(16) => n50, A(15) => n48, A(14) => n45, A(13) => 
                           n43, A(12) => n41, A(11) => n39, A(10) => n37, A(9) 
                           => n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) 
                           => n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) 
                           => n19, A(0) => n17, p(32) => q_0_1_42_port, p(31) 
                           => q_0_1_41_port, p(30) => q_0_2_40_port, p(29) => 
                           q_0_2_39_port, p(28) => q_0_3_38_port, p(27) => 
                           q_0_3_37_port, p(26) => q_0_4_36_port, p(25) => 
                           q_0_5_35_port, p(24) => q_0_5_34_port, p(23) => 
                           q_0_5_33_port, p(22) => q_0_5_32_port, p(21) => 
                           q_0_5_31_port, p(20) => q_0_5_30_port, p(19) => 
                           q_0_5_29_port, p(18) => q_0_5_28_port, p(17) => 
                           q_0_5_27_port, p(16) => q_0_5_26_port, p(15) => 
                           q_0_5_25_port, p(14) => q_0_5_24_port, p(13) => 
                           q_0_5_23_port, p(12) => q_0_5_22_port, p(11) => 
                           q_0_5_21_port, p(10) => q_0_5_20_port, p(9) => 
                           q_0_5_19_port, p(8) => q_0_5_18_port, p(7) => 
                           q_0_5_17_port, p(6) => q_0_5_16_port, p(5) => 
                           q_0_5_15_port, p(4) => q_0_5_14_port, p(3) => 
                           q_0_5_13_port, p(2) => q_0_5_12_port, p(1) => 
                           q_0_5_11_port, p(0) => q_0_5_10_port);
   encI_7 : ENC_11 port map( b(2) => B(13), b(1) => B(12), b(0) => B(11), A(31)
                           => n79, A(30) => n77, A(29) => n75, A(28) => n73, 
                           A(27) => n71, A(26) => n69, A(25) => n67, A(24) => 
                           n65, A(23) => n63, A(22) => n61, A(21) => n60, A(20)
                           => n57, A(19) => n55, A(18) => n53, A(17) => n51, 
                           A(16) => n49, A(15) => n47, A(14) => n45, A(13) => 
                           n43, A(12) => n41, A(11) => n39, A(10) => n37, A(9) 
                           => n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) 
                           => n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) 
                           => n19, A(0) => n17, p(32) => q_0_1_44_port, p(31) 
                           => q_0_1_43_port, p(30) => q_0_2_42_port, p(29) => 
                           q_0_2_41_port, p(28) => q_0_3_40_port, p(27) => 
                           q_0_3_39_port, p(26) => q_0_4_38_port, p(25) => 
                           q_0_4_37_port, p(24) => q_0_5_36_port, p(23) => 
                           q_0_6_35_port, p(22) => q_0_6_34_port, p(21) => 
                           q_0_6_33_port, p(20) => q_0_6_32_port, p(19) => 
                           q_0_6_31_port, p(18) => q_0_6_30_port, p(17) => 
                           q_0_6_29_port, p(16) => q_0_6_28_port, p(15) => 
                           q_0_6_27_port, p(14) => q_0_6_26_port, p(13) => 
                           q_0_6_25_port, p(12) => q_0_6_24_port, p(11) => 
                           q_0_6_23_port, p(10) => q_0_6_22_port, p(9) => 
                           q_0_6_21_port, p(8) => q_0_6_20_port, p(7) => 
                           q_0_6_19_port, p(6) => q_0_6_18_port, p(5) => 
                           q_0_6_17_port, p(4) => q_0_6_16_port, p(3) => 
                           q_0_6_15_port, p(2) => q_0_6_14_port, p(1) => 
                           q_0_6_13_port, p(0) => q_0_6_12_port);
   encI_8 : ENC_10 port map( b(2) => B(15), b(1) => B(14), b(0) => B(13), A(31)
                           => n79, A(30) => n77, A(29) => n75, A(28) => n73, 
                           A(27) => n71, A(26) => n69, A(25) => n67, A(24) => 
                           n65, A(23) => n63, A(22) => n61, A(21) => n59, A(20)
                           => n57, A(19) => n55, A(18) => n53, A(17) => n51, 
                           A(16) => n49, A(15) => n47, A(14) => n45, A(13) => 
                           n43, A(12) => n41, A(11) => n39, A(10) => n37, A(9) 
                           => n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) 
                           => n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) 
                           => n19, A(0) => n17, p(32) => q_0_1_46_port, p(31) 
                           => q_0_1_45_port, p(30) => q_0_2_44_port, p(29) => 
                           q_0_2_43_port, p(28) => q_0_3_42_port, p(27) => 
                           q_0_3_41_port, p(26) => q_0_4_40_port, p(25) => 
                           q_0_4_39_port, p(24) => q_0_5_38_port, p(23) => 
                           q_0_5_37_port, p(22) => q_0_6_36_port, p(21) => 
                           q_0_7_35_port, p(20) => q_0_7_34_port, p(19) => 
                           q_0_7_33_port, p(18) => q_0_7_32_port, p(17) => 
                           q_0_7_31_port, p(16) => q_0_7_30_port, p(15) => 
                           q_0_7_29_port, p(14) => q_0_7_28_port, p(13) => 
                           q_0_7_27_port, p(12) => q_0_7_26_port, p(11) => 
                           q_0_7_25_port, p(10) => q_0_7_24_port, p(9) => 
                           q_0_7_23_port, p(8) => q_0_7_22_port, p(7) => 
                           q_0_7_21_port, p(6) => q_0_7_20_port, p(5) => 
                           q_0_7_19_port, p(4) => q_0_7_18_port, p(3) => 
                           q_0_7_17_port, p(2) => q_0_7_16_port, p(1) => 
                           q_0_7_15_port, p(0) => q_0_7_14_port);
   encI_9 : ENC_9 port map( b(2) => B(17), b(1) => B(16), b(0) => B(15), A(31) 
                           => n80, A(30) => n77, A(29) => n75, A(28) => n73, 
                           A(27) => n71, A(26) => n69, A(25) => n67, A(24) => 
                           n65, A(23) => n63, A(22) => n61, A(21) => n59, A(20)
                           => n57, A(19) => n55, A(18) => n53, A(17) => n51, 
                           A(16) => n49, A(15) => n47, A(14) => n45, A(13) => 
                           n43, A(12) => n41, A(11) => n39, A(10) => n37, A(9) 
                           => n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) 
                           => n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) 
                           => n19, A(0) => n17, p(32) => q_0_1_48_port, p(31) 
                           => q_0_1_47_port, p(30) => q_0_2_46_port, p(29) => 
                           q_0_2_45_port, p(28) => q_0_3_44_port, p(27) => 
                           q_0_3_43_port, p(26) => q_0_4_42_port, p(25) => 
                           q_0_4_41_port, p(24) => q_0_5_40_port, p(23) => 
                           q_0_5_39_port, p(22) => q_0_6_38_port, p(21) => 
                           q_0_6_37_port, p(20) => q_0_7_36_port, p(19) => 
                           q_0_8_35_port, p(18) => q_0_8_34_port, p(17) => 
                           q_0_8_33_port, p(16) => q_0_8_32_port, p(15) => 
                           q_0_8_31_port, p(14) => q_0_8_30_port, p(13) => 
                           q_0_8_29_port, p(12) => q_0_8_28_port, p(11) => 
                           q_0_8_27_port, p(10) => q_0_8_26_port, p(9) => 
                           q_0_8_25_port, p(8) => q_0_8_24_port, p(7) => 
                           q_0_8_23_port, p(6) => q_0_8_22_port, p(5) => 
                           q_0_8_21_port, p(4) => q_0_8_20_port, p(3) => 
                           q_0_8_19_port, p(2) => q_0_8_18_port, p(1) => 
                           q_0_8_17_port, p(0) => q_0_8_16_port);
   encI_10 : ENC_8 port map( b(2) => B(19), b(1) => B(18), b(0) => B(17), A(31)
                           => n80, A(30) => n77, A(29) => n75, A(28) => n73, 
                           A(27) => n71, A(26) => n69, A(25) => n67, A(24) => 
                           n65, A(23) => n63, A(22) => n61, A(21) => n59, A(20)
                           => n57, A(19) => n55, A(18) => n53, A(17) => n51, 
                           A(16) => n49, A(15) => n47, A(14) => n45, A(13) => 
                           n43, A(12) => n41, A(11) => n39, A(10) => n37, A(9) 
                           => n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) 
                           => n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) 
                           => n19, A(0) => n17, p(32) => q_0_1_50_port, p(31) 
                           => q_0_1_49_port, p(30) => q_0_2_48_port, p(29) => 
                           q_0_2_47_port, p(28) => q_0_3_46_port, p(27) => 
                           q_0_3_45_port, p(26) => q_0_4_44_port, p(25) => 
                           q_0_4_43_port, p(24) => q_0_5_42_port, p(23) => 
                           q_0_5_41_port, p(22) => q_0_6_40_port, p(21) => 
                           q_0_6_39_port, p(20) => q_0_7_38_port, p(19) => 
                           q_0_7_37_port, p(18) => q_0_8_36_port, p(17) => 
                           q_0_9_35_port, p(16) => q_0_9_34_port, p(15) => 
                           q_0_9_33_port, p(14) => q_0_9_32_port, p(13) => 
                           q_0_9_31_port, p(12) => q_0_9_30_port, p(11) => 
                           q_0_9_29_port, p(10) => q_0_9_28_port, p(9) => 
                           q_0_9_27_port, p(8) => q_0_9_26_port, p(7) => 
                           q_0_9_25_port, p(6) => q_0_9_24_port, p(5) => 
                           q_0_9_23_port, p(4) => q_0_9_22_port, p(3) => 
                           q_0_9_21_port, p(2) => q_0_9_20_port, p(1) => 
                           q_0_9_19_port, p(0) => q_0_9_18_port);
   encI_11 : ENC_7 port map( b(2) => B(21), b(1) => B(20), b(0) => B(19), A(31)
                           => n80, A(30) => n78, A(29) => n76, A(28) => n73, 
                           A(27) => n71, A(26) => n69, A(25) => n67, A(24) => 
                           n65, A(23) => n63, A(22) => n61, A(21) => n59, A(20)
                           => n57, A(19) => n55, A(18) => n53, A(17) => n51, 
                           A(16) => n49, A(15) => n47, A(14) => n45, A(13) => 
                           n43, A(12) => n41, A(11) => n39, A(10) => n37, A(9) 
                           => n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) 
                           => n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) 
                           => n19, A(0) => n17, p(32) => q_0_1_52_port, p(31) 
                           => q_0_1_51_port, p(30) => q_0_2_50_port, p(29) => 
                           q_0_2_49_port, p(28) => q_0_3_48_port, p(27) => 
                           q_0_3_47_port, p(26) => q_0_4_46_port, p(25) => 
                           q_0_4_45_port, p(24) => q_0_5_44_port, p(23) => 
                           q_0_5_43_port, p(22) => q_0_6_42_port, p(21) => 
                           q_0_6_41_port, p(20) => q_0_7_40_port, p(19) => 
                           q_0_7_39_port, p(18) => q_0_8_38_port, p(17) => 
                           q_0_8_37_port, p(16) => q_0_9_36_port, p(15) => 
                           q_0_10_35_port, p(14) => q_0_10_34_port, p(13) => 
                           q_0_10_33_port, p(12) => q_0_10_32_port, p(11) => 
                           q_0_10_31_port, p(10) => q_0_10_30_port, p(9) => 
                           q_0_10_29_port, p(8) => q_0_10_28_port, p(7) => 
                           q_0_10_27_port, p(6) => q_0_10_26_port, p(5) => 
                           q_0_10_25_port, p(4) => q_0_10_24_port, p(3) => 
                           q_0_10_23_port, p(2) => q_0_10_22_port, p(1) => 
                           q_0_10_21_port, p(0) => q_0_10_20_port);
   encI_12 : ENC_6 port map( b(2) => n3, b(1) => B(22), b(0) => B(21), A(31) =>
                           n80, A(30) => n78, A(29) => n76, A(28) => n73, A(27)
                           => n71, A(26) => n69, A(25) => n67, A(24) => n65, 
                           A(23) => n63, A(22) => n61, A(21) => n59, A(20) => 
                           n57, A(19) => n55, A(18) => n53, A(17) => n51, A(16)
                           => n49, A(15) => n47, A(14) => n45, A(13) => n43, 
                           A(12) => n41, A(11) => n39, A(10) => n37, A(9) => 
                           n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) => 
                           n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) => 
                           n19, A(0) => n17, p(32) => q_0_1_54_port, p(31) => 
                           q_0_1_53_port, p(30) => q_0_2_52_port, p(29) => 
                           q_0_2_51_port, p(28) => q_0_3_50_port, p(27) => 
                           q_0_3_49_port, p(26) => q_0_4_48_port, p(25) => 
                           q_0_4_47_port, p(24) => q_0_5_46_port, p(23) => 
                           q_0_5_45_port, p(22) => q_0_6_44_port, p(21) => 
                           q_0_6_43_port, p(20) => q_0_7_42_port, p(19) => 
                           q_0_7_41_port, p(18) => q_0_8_40_port, p(17) => 
                           q_0_8_39_port, p(16) => q_0_9_38_port, p(15) => 
                           q_0_9_37_port, p(14) => q_0_10_36_port, p(13) => 
                           q_0_11_35_port, p(12) => q_0_11_34_port, p(11) => 
                           q_0_11_33_port, p(10) => q_0_11_32_port, p(9) => 
                           q_0_11_31_port, p(8) => q_0_11_30_port, p(7) => 
                           q_0_11_29_port, p(6) => q_0_11_28_port, p(5) => 
                           q_0_11_27_port, p(4) => q_0_11_26_port, p(3) => 
                           q_0_11_25_port, p(2) => q_0_11_24_port, p(1) => 
                           q_0_11_23_port, p(0) => q_0_11_22_port);
   encI_13 : ENC_5 port map( b(2) => B(25), b(1) => B(24), b(0) => B(23), A(31)
                           => n80, A(30) => n78, A(29) => n76, A(28) => n74, 
                           A(27) => n72, A(26) => n70, A(25) => n68, A(24) => 
                           n66, A(23) => n64, A(22) => n61, A(21) => n59, A(20)
                           => n57, A(19) => n55, A(18) => n53, A(17) => n51, 
                           A(16) => n49, A(15) => n47, A(14) => n45, A(13) => 
                           n43, A(12) => n41, A(11) => n39, A(10) => n37, A(9) 
                           => n35, A(8) => n33, A(7) => n31, A(6) => n29, A(5) 
                           => n27, A(4) => n25, A(3) => n23, A(2) => n21, A(1) 
                           => n19, A(0) => n17, p(32) => q_0_1_56_port, p(31) 
                           => q_0_1_55_port, p(30) => q_0_2_54_port, p(29) => 
                           q_0_2_53_port, p(28) => q_0_3_52_port, p(27) => 
                           q_0_3_51_port, p(26) => q_0_4_50_port, p(25) => 
                           q_0_4_49_port, p(24) => q_0_5_48_port, p(23) => 
                           q_0_5_47_port, p(22) => q_0_6_46_port, p(21) => 
                           q_0_6_45_port, p(20) => q_0_7_44_port, p(19) => 
                           q_0_7_43_port, p(18) => q_0_8_42_port, p(17) => 
                           q_0_8_41_port, p(16) => q_0_9_40_port, p(15) => 
                           q_0_9_39_port, p(14) => q_0_10_38_port, p(13) => 
                           q_0_10_37_port, p(12) => q_0_11_36_port, p(11) => 
                           q_0_12_35_port, p(10) => q_0_12_34_port, p(9) => 
                           q_0_12_33_port, p(8) => q_0_12_32_port, p(7) => 
                           q_0_12_31_port, p(6) => q_0_12_30_port, p(5) => 
                           q_0_12_29_port, p(4) => q_0_12_28_port, p(3) => 
                           q_0_12_27_port, p(2) => q_0_12_26_port, p(1) => 
                           q_0_12_25_port, p(0) => q_0_12_24_port);
   encI_14 : ENC_4 port map( b(2) => B(27), b(1) => B(26), b(0) => B(25), A(31)
                           => n80, A(30) => n78, A(29) => n76, A(28) => n74, 
                           A(27) => n72, A(26) => n70, A(25) => n68, A(24) => 
                           n66, A(23) => n64, A(22) => n62, A(21) => n60, A(20)
                           => n57, A(19) => n55, A(18) => n53, A(17) => n51, 
                           A(16) => n49, A(15) => n47, A(14) => n46, A(13) => 
                           n44, A(12) => n42, A(11) => n40, A(10) => n38, A(9) 
                           => n36, A(8) => n34, A(7) => n32, A(6) => n30, A(5) 
                           => n28, A(4) => n26, A(3) => n24, A(2) => n22, A(1) 
                           => n20, A(0) => n18, p(32) => q_0_1_58_port, p(31) 
                           => q_0_1_57_port, p(30) => q_0_2_56_port, p(29) => 
                           q_0_2_55_port, p(28) => q_0_3_54_port, p(27) => 
                           q_0_3_53_port, p(26) => q_0_4_52_port, p(25) => 
                           q_0_4_51_port, p(24) => q_0_5_50_port, p(23) => 
                           q_0_5_49_port, p(22) => q_0_6_48_port, p(21) => 
                           q_0_6_47_port, p(20) => q_0_7_46_port, p(19) => 
                           q_0_7_45_port, p(18) => q_0_8_44_port, p(17) => 
                           q_0_8_43_port, p(16) => q_0_9_42_port, p(15) => 
                           q_0_9_41_port, p(14) => q_0_10_40_port, p(13) => 
                           q_0_10_39_port, p(12) => q_0_11_38_port, p(11) => 
                           q_0_11_37_port, p(10) => q_0_12_36_port, p(9) => 
                           q_0_13_35_port, p(8) => q_0_13_34_port, p(7) => 
                           q_0_13_33_port, p(6) => q_0_13_32_port, p(5) => 
                           q_0_13_31_port, p(4) => q_0_13_30_port, p(3) => 
                           q_0_13_29_port, p(2) => q_0_13_28_port, p(1) => 
                           q_0_13_27_port, p(0) => q_0_13_26_port);
   encI_15 : ENC_3 port map( b(2) => B(29), b(1) => B(28), b(0) => B(27), A(31)
                           => n80, A(30) => n77, A(29) => n75, A(28) => n74, 
                           A(27) => n72, A(26) => n70, A(25) => n68, A(24) => 
                           n66, A(23) => n64, A(22) => n62, A(21) => n60, A(20)
                           => n58, A(19) => n56, A(18) => n53, A(17) => n51, 
                           A(16) => n49, A(15) => n47, A(14) => n46, A(13) => 
                           n44, A(12) => n42, A(11) => n40, A(10) => n38, A(9) 
                           => n36, A(8) => n34, A(7) => n32, A(6) => n30, A(5) 
                           => n28, A(4) => n26, A(3) => n24, A(2) => n22, A(1) 
                           => n20, A(0) => n18, p(32) => q_0_1_60_port, p(31) 
                           => q_0_1_59_port, p(30) => q_0_2_58_port, p(29) => 
                           q_0_2_57_port, p(28) => q_0_3_56_port, p(27) => 
                           q_0_3_55_port, p(26) => q_0_4_54_port, p(25) => 
                           q_0_4_53_port, p(24) => q_0_5_52_port, p(23) => 
                           q_0_5_51_port, p(22) => q_0_6_50_port, p(21) => 
                           q_0_6_49_port, p(20) => q_0_7_48_port, p(19) => 
                           q_0_7_47_port, p(18) => q_0_8_46_port, p(17) => 
                           q_0_8_45_port, p(16) => q_0_9_44_port, p(15) => 
                           q_0_9_43_port, p(14) => q_0_10_42_port, p(13) => 
                           q_0_10_41_port, p(12) => q_0_11_40_port, p(11) => 
                           q_0_11_39_port, p(10) => q_0_12_38_port, p(9) => 
                           q_0_12_37_port, p(8) => q_0_13_36_port, p(7) => 
                           q_0_14_35_port, p(6) => q_0_14_34_port, p(5) => 
                           q_0_14_33_port, p(4) => q_0_14_32_port, p(3) => 
                           q_0_14_31_port, p(2) => q_0_14_30_port, p(1) => 
                           q_0_14_29_port, p(0) => q_0_14_28_port);
   encI_16 : ENC_2 port map( b(2) => B(31), b(1) => B(30), b(0) => B(29), A(31)
                           => n80, A(30) => n78, A(29) => n76, A(28) => n74, 
                           A(27) => n72, A(26) => n70, A(25) => n68, A(24) => 
                           n66, A(23) => n64, A(22) => n62, A(21) => n60, A(20)
                           => n58, A(19) => n56, A(18) => n54, A(17) => n52, 
                           A(16) => n49, A(15) => n47, A(14) => n46, A(13) => 
                           n44, A(12) => n42, A(11) => n40, A(10) => n38, A(9) 
                           => n36, A(8) => n34, A(7) => n32, A(6) => n30, A(5) 
                           => n28, A(4) => n26, A(3) => n24, A(2) => n22, A(1) 
                           => n20, A(0) => n18, p(32) => q_0_1_62_port, p(31) 
                           => q_0_1_61_port, p(30) => q_0_2_60_port, p(29) => 
                           q_0_2_59_port, p(28) => q_0_3_58_port, p(27) => 
                           q_0_3_57_port, p(26) => q_0_4_56_port, p(25) => 
                           q_0_4_55_port, p(24) => q_0_5_54_port, p(23) => 
                           q_0_5_53_port, p(22) => q_0_6_52_port, p(21) => 
                           q_0_6_51_port, p(20) => q_0_7_50_port, p(19) => 
                           q_0_7_49_port, p(18) => q_0_8_48_port, p(17) => 
                           q_0_8_47_port, p(16) => q_0_9_46_port, p(15) => 
                           q_0_9_45_port, p(14) => q_0_10_44_port, p(13) => 
                           q_0_10_43_port, p(12) => q_0_11_42_port, p(11) => 
                           q_0_11_41_port, p(10) => q_0_12_40_port, p(9) => 
                           q_0_12_39_port, p(8) => q_0_13_38_port, p(7) => 
                           q_0_13_37_port, p(6) => q_0_14_36_port, p(5) => 
                           q_0_15_35_port, p(4) => q_0_15_34_port, p(3) => 
                           q_0_15_33_port, p(2) => q_0_15_32_port, p(1) => 
                           q_0_15_31_port, p(0) => q_0_15_30_port);
   encI_17 : ENC_1 port map( b(2) => X_Logic0_port, b(1) => X_Logic0_port, b(0)
                           => B(31), A(31) => n80, A(30) => n77, A(29) => n75, 
                           A(28) => n74, A(27) => n72, A(26) => n70, A(25) => 
                           n68, A(24) => n66, A(23) => n64, A(22) => n62, A(21)
                           => n60, A(20) => n58, A(19) => n56, A(18) => n54, 
                           A(17) => n52, A(16) => n50, A(15) => n48, A(14) => 
                           n46, A(13) => n44, A(12) => n42, A(11) => n40, A(10)
                           => n38, A(9) => n36, A(8) => n34, A(7) => n32, A(6) 
                           => n30, A(5) => n28, A(4) => n26, A(3) => n24, A(2) 
                           => n22, A(1) => n20, A(0) => n18, p(32) => n_1042, 
                           p(31) => q_0_1_63_port, p(30) => q_0_2_62_port, 
                           p(29) => q_0_2_61_port, p(28) => q_0_3_60_port, 
                           p(27) => q_0_3_59_port, p(26) => q_0_4_58_port, 
                           p(25) => q_0_4_57_port, p(24) => q_0_5_56_port, 
                           p(23) => q_0_5_55_port, p(22) => q_0_6_54_port, 
                           p(21) => q_0_6_53_port, p(20) => q_0_7_52_port, 
                           p(19) => q_0_7_51_port, p(18) => q_0_8_50_port, 
                           p(17) => q_0_8_49_port, p(16) => q_0_9_48_port, 
                           p(15) => q_0_9_47_port, p(14) => q_0_10_46_port, 
                           p(13) => q_0_10_45_port, p(12) => q_0_11_44_port, 
                           p(11) => q_0_11_43_port, p(10) => q_0_12_42_port, 
                           p(9) => q_0_12_41_port, p(8) => q_0_13_40_port, p(7)
                           => q_0_13_39_port, p(6) => q_0_14_38_port, p(5) => 
                           q_0_14_37_port, p(4) => q_0_15_36_port, p(3) => 
                           q_0_16_35_port, p(2) => q_0_16_34_port, p(1) => 
                           q_0_16_33_port, p(0) => q_0_16_32_port);
   HA_R_0_0_24 : HA_0 port map( A => q_0_0_24_port, B => q_0_1_24_port, S => 
                           q_1_0_24_port, C => q_1_1_25_port);
   HA_R_0_0_25 : HA_43 port map( A => q_0_0_25_port, B => q_0_1_25_port, S => 
                           q_1_0_25_port, C => q_1_1_26_port);
   FA_C_0_0_26 : FA_0 port map( A => q_0_0_26_port, B => q_0_1_26_port, Ci => 
                           q_0_2_26_port, S => q_1_0_26_port, Co => 
                           q_1_1_27_port);
   FA_C_0_0_27 : FA_607 port map( A => q_0_0_27_port, B => q_0_1_27_port, Ci =>
                           q_0_2_27_port, S => q_1_0_27_port, Co => 
                           q_1_1_28_port);
   FA_C_0_0_28 : FA_606 port map( A => q_0_0_28_port, B => q_0_1_28_port, Ci =>
                           q_0_2_28_port, S => q_1_0_28_port, Co => 
                           q_1_1_29_port);
   FA_C_0_0_29 : FA_605 port map( A => q_0_0_29_port, B => q_0_1_29_port, Ci =>
                           q_0_2_29_port, S => q_1_0_29_port, Co => 
                           q_1_1_30_port);
   FA_C_0_0_30 : FA_604 port map( A => q_0_0_30_port, B => q_0_1_30_port, Ci =>
                           q_0_2_30_port, S => q_1_0_30_port, Co => 
                           q_1_1_31_port);
   FA_C_0_0_31 : FA_603 port map( A => q_0_0_31_port, B => q_0_1_31_port, Ci =>
                           q_0_2_31_port, S => q_1_0_31_port, Co => 
                           q_1_1_32_port);
   FA_C_0_0_32 : FA_602 port map( A => q_0_0_32_port, B => q_0_1_32_port, Ci =>
                           q_0_2_32_port, S => q_1_0_32_port, Co => 
                           q_1_1_33_port);
   FA_C_0_0_33 : FA_601 port map( A => n15, B => q_0_1_33_port, Ci => 
                           q_0_2_33_port, S => q_1_0_33_port, Co => 
                           q_1_1_34_port);
   FA_C_0_0_34 : FA_600 port map( A => n12, B => q_0_1_34_port, Ci => 
                           q_0_2_34_port, S => q_1_0_34_port, Co => 
                           q_1_1_35_port);
   FA_C_0_0_35 : FA_599 port map( A => n96, B => n95, Ci => q_0_2_35_port, S =>
                           q_1_0_35_port, Co => q_1_1_36_port);
   FA_C_0_0_36 : FA_598 port map( A => X_Logic1_port, B => q_0_1_36_port, Ci =>
                           q_0_2_36_port, S => q_1_0_36_port, Co => 
                           q_1_1_37_port);
   FA_C_0_0_37 : FA_597 port map( A => n94, B => q_0_1_37_port, Ci => 
                           q_0_2_37_port, S => q_1_0_37_port, Co => 
                           q_1_1_38_port);
   FA_C_0_0_38 : FA_596 port map( A => X_Logic1_port, B => q_0_1_38_port, Ci =>
                           q_0_2_38_port, S => q_1_0_38_port, Co => 
                           q_1_1_39_port);
   FA_C_0_0_39 : FA_595 port map( A => n93, B => q_0_1_39_port, Ci => 
                           q_0_2_39_port, S => q_1_0_39_port, Co => 
                           q_1_1_40_port);
   FA_C_0_0_40 : FA_594 port map( A => X_Logic1_port, B => q_0_1_40_port, Ci =>
                           q_0_2_40_port, S => q_1_0_40_port, Co => 
                           q_1_1_41_port);
   FA_C_0_0_41 : FA_593 port map( A => n92, B => q_0_1_41_port, Ci => 
                           q_0_2_41_port, S => q_1_0_41_port, Co => 
                           q_1_1_42_port);
   HA_L_0_0_42 : HA_42 port map( A => X_Logic1_port, B => q_0_1_42_port, S => 
                           q_1_0_42_port, C => q_1_0_43_port);
   HA_R_0_3_26 : HA_41 port map( A => q_0_3_26_port, B => q_0_4_26_port, S => 
                           q_1_2_26_port, C => q_1_3_27_port);
   HA_R_0_3_27 : HA_40 port map( A => q_0_3_27_port, B => q_0_4_27_port, S => 
                           q_1_2_27_port, C => q_1_3_28_port);
   FA_C_0_3_28 : FA_592 port map( A => q_0_3_28_port, B => q_0_4_28_port, Ci =>
                           q_0_5_28_port, S => q_1_2_28_port, Co => 
                           q_1_3_29_port);
   FA_C_0_3_29 : FA_591 port map( A => q_0_3_29_port, B => q_0_4_29_port, Ci =>
                           q_0_5_29_port, S => q_1_2_29_port, Co => 
                           q_1_3_30_port);
   FA_C_0_3_30 : FA_590 port map( A => q_0_3_30_port, B => q_0_4_30_port, Ci =>
                           q_0_5_30_port, S => q_1_2_30_port, Co => 
                           q_1_3_31_port);
   FA_C_0_3_31 : FA_589 port map( A => q_0_3_31_port, B => q_0_4_31_port, Ci =>
                           q_0_5_31_port, S => q_1_2_31_port, Co => 
                           q_1_3_32_port);
   FA_C_0_3_32 : FA_588 port map( A => q_0_3_32_port, B => q_0_4_32_port, Ci =>
                           q_0_5_32_port, S => q_1_2_32_port, Co => 
                           q_1_3_33_port);
   FA_C_0_3_33 : FA_587 port map( A => q_0_3_33_port, B => q_0_4_33_port, Ci =>
                           q_0_5_33_port, S => q_1_2_33_port, Co => 
                           q_1_3_34_port);
   FA_C_0_3_34 : FA_586 port map( A => q_0_3_34_port, B => q_0_4_34_port, Ci =>
                           q_0_5_34_port, S => q_1_2_34_port, Co => 
                           q_1_3_35_port);
   FA_C_0_3_35 : FA_585 port map( A => q_0_3_35_port, B => q_0_4_35_port, Ci =>
                           q_0_5_35_port, S => q_1_2_35_port, Co => 
                           q_1_3_36_port);
   FA_C_0_3_36 : FA_584 port map( A => q_0_3_36_port, B => q_0_4_36_port, Ci =>
                           q_0_5_36_port, S => q_1_2_36_port, Co => 
                           q_1_3_37_port);
   FA_C_0_3_37 : FA_583 port map( A => q_0_3_37_port, B => q_0_4_37_port, Ci =>
                           q_0_5_37_port, S => q_1_2_37_port, Co => 
                           q_1_3_38_port);
   FA_C_0_3_38 : FA_582 port map( A => q_0_3_38_port, B => q_0_4_38_port, Ci =>
                           q_0_5_38_port, S => q_1_2_38_port, Co => 
                           q_1_3_39_port);
   FA_C_0_3_39 : FA_581 port map( A => q_0_3_39_port, B => q_0_4_39_port, Ci =>
                           q_0_5_39_port, S => q_1_2_39_port, Co => 
                           q_1_3_40_port);
   HA_L_0_3_40 : HA_39 port map( A => q_0_3_40_port, B => q_0_4_40_port, S => 
                           q_1_2_40_port, C => q_1_2_41_port);
   HA_R_0_6_28 : HA_38 port map( A => q_0_6_28_port, B => q_0_7_28_port, S => 
                           q_1_4_28_port, C => q_1_5_29_port);
   HA_R_0_6_29 : HA_37 port map( A => q_0_6_29_port, B => q_0_7_29_port, S => 
                           q_1_4_29_port, C => q_1_5_30_port);
   FA_C_0_6_30 : FA_580 port map( A => q_0_6_30_port, B => q_0_7_30_port, Ci =>
                           q_0_8_30_port, S => q_1_4_30_port, Co => 
                           q_1_5_31_port);
   FA_C_0_6_31 : FA_579 port map( A => q_0_6_31_port, B => q_0_7_31_port, Ci =>
                           q_0_8_31_port, S => q_1_4_31_port, Co => 
                           q_1_5_32_port);
   FA_C_0_6_32 : FA_578 port map( A => q_0_6_32_port, B => q_0_7_32_port, Ci =>
                           q_0_8_32_port, S => q_1_4_32_port, Co => 
                           q_1_5_33_port);
   FA_C_0_6_33 : FA_577 port map( A => q_0_6_33_port, B => q_0_7_33_port, Ci =>
                           q_0_8_33_port, S => q_1_4_33_port, Co => 
                           q_1_5_34_port);
   FA_C_0_6_34 : FA_576 port map( A => q_0_6_34_port, B => q_0_7_34_port, Ci =>
                           q_0_8_34_port, S => q_1_4_34_port, Co => 
                           q_1_5_35_port);
   FA_C_0_6_35 : FA_575 port map( A => q_0_6_35_port, B => q_0_7_35_port, Ci =>
                           q_0_8_35_port, S => q_1_4_35_port, Co => 
                           q_1_5_36_port);
   FA_C_0_6_36 : FA_574 port map( A => q_0_6_36_port, B => q_0_7_36_port, Ci =>
                           q_0_8_36_port, S => q_1_4_36_port, Co => 
                           q_1_5_37_port);
   FA_C_0_6_37 : FA_573 port map( A => q_0_6_37_port, B => q_0_7_37_port, Ci =>
                           q_0_8_37_port, S => q_1_4_37_port, Co => 
                           q_1_5_38_port);
   HA_L_0_6_38 : HA_36 port map( A => q_0_6_38_port, B => q_0_7_38_port, S => 
                           q_1_4_38_port, C => q_1_4_39_port);
   HA_R_0_9_30 : HA_35 port map( A => q_0_9_30_port, B => q_0_10_30_port, S => 
                           q_1_6_30_port, C => q_1_7_31_port);
   HA_R_0_9_31 : HA_34 port map( A => q_0_9_31_port, B => q_0_10_31_port, S => 
                           q_1_6_31_port, C => q_1_7_32_port);
   FA_C_0_9_32 : FA_572 port map( A => q_0_9_32_port, B => q_0_10_32_port, Ci 
                           => q_0_11_32_port, S => q_1_6_32_port, Co => 
                           q_1_7_33_port);
   FA_C_0_9_33 : FA_571 port map( A => q_0_9_33_port, B => q_0_10_33_port, Ci 
                           => q_0_11_33_port, S => q_1_6_33_port, Co => 
                           q_1_7_34_port);
   FA_C_0_9_34 : FA_570 port map( A => q_0_9_34_port, B => q_0_10_34_port, Ci 
                           => q_0_11_34_port, S => q_1_6_34_port, Co => 
                           q_1_7_35_port);
   FA_C_0_9_35 : FA_569 port map( A => q_0_9_35_port, B => q_0_10_35_port, Ci 
                           => q_0_11_35_port, S => q_1_6_35_port, Co => 
                           q_1_7_36_port);
   HA_L_0_9_36 : HA_33 port map( A => q_0_9_36_port, B => q_0_10_36_port, S => 
                           q_1_6_36_port, C => q_1_6_37_port);
   HA_R_1_0_16 : HA_32 port map( A => q_0_0_16_port, B => q_0_1_16_port, S => 
                           q_2_0_16_port, C => q_2_1_17_port);
   HA_R_1_0_17 : HA_31 port map( A => q_0_0_17_port, B => q_0_1_17_port, S => 
                           q_2_0_17_port, C => q_2_1_18_port);
   FA_C_1_0_18 : FA_568 port map( A => q_0_0_18_port, B => q_0_1_18_port, Ci =>
                           q_0_2_18_port, S => q_2_0_18_port, Co => 
                           q_2_1_19_port);
   FA_C_1_0_19 : FA_567 port map( A => q_0_0_19_port, B => q_0_1_19_port, Ci =>
                           q_0_2_19_port, S => q_2_0_19_port, Co => 
                           q_2_1_20_port);
   FA_C_1_0_20 : FA_566 port map( A => q_0_0_20_port, B => q_0_1_20_port, Ci =>
                           q_0_2_20_port, S => q_2_0_20_port, Co => 
                           q_2_1_21_port);
   FA_C_1_0_21 : FA_565 port map( A => q_0_0_21_port, B => q_0_1_21_port, Ci =>
                           q_0_2_21_port, S => q_2_0_21_port, Co => 
                           q_2_1_22_port);
   FA_C_1_0_22 : FA_564 port map( A => q_0_0_22_port, B => q_0_1_22_port, Ci =>
                           q_0_2_22_port, S => q_2_0_22_port, Co => 
                           q_2_1_23_port);
   FA_C_1_0_23 : FA_563 port map( A => q_0_0_23_port, B => q_0_1_23_port, Ci =>
                           q_0_2_23_port, S => q_2_0_23_port, Co => 
                           q_2_1_24_port);
   FA_C_1_0_24 : FA_562 port map( A => q_1_0_24_port, B => q_0_2_24_port, Ci =>
                           q_0_3_24_port, S => q_2_0_24_port, Co => 
                           q_2_1_25_port);
   FA_C_1_0_25 : FA_561 port map( A => q_1_0_25_port, B => q_1_1_25_port, Ci =>
                           q_0_2_25_port, S => q_2_0_25_port, Co => 
                           q_2_1_26_port);
   FA_C_1_0_26 : FA_560 port map( A => q_1_0_26_port, B => q_1_1_26_port, Ci =>
                           q_1_2_26_port, S => q_2_0_26_port, Co => 
                           q_2_1_27_port);
   FA_C_1_0_27 : FA_559 port map( A => q_1_0_27_port, B => q_1_1_27_port, Ci =>
                           q_1_2_27_port, S => q_2_0_27_port, Co => 
                           q_2_1_28_port);
   FA_C_1_0_28 : FA_558 port map( A => q_1_0_28_port, B => q_1_1_28_port, Ci =>
                           q_1_2_28_port, S => q_2_0_28_port, Co => 
                           q_2_1_29_port);
   FA_C_1_0_29 : FA_557 port map( A => q_1_0_29_port, B => q_1_1_29_port, Ci =>
                           q_1_2_29_port, S => q_2_0_29_port, Co => 
                           q_2_1_30_port);
   FA_C_1_0_30 : FA_556 port map( A => q_1_0_30_port, B => q_1_1_30_port, Ci =>
                           q_1_2_30_port, S => q_2_0_30_port, Co => 
                           q_2_1_31_port);
   FA_C_1_0_31 : FA_555 port map( A => q_1_0_31_port, B => q_1_1_31_port, Ci =>
                           q_1_2_31_port, S => q_2_0_31_port, Co => 
                           q_2_1_32_port);
   FA_C_1_0_32 : FA_554 port map( A => q_1_0_32_port, B => q_1_1_32_port, Ci =>
                           q_1_2_32_port, S => q_2_0_32_port, Co => 
                           q_2_1_33_port);
   FA_C_1_0_33 : FA_553 port map( A => q_1_0_33_port, B => q_1_1_33_port, Ci =>
                           q_1_2_33_port, S => q_2_0_33_port, Co => 
                           q_2_1_34_port);
   FA_C_1_0_34 : FA_552 port map( A => q_1_0_34_port, B => q_1_1_34_port, Ci =>
                           q_1_2_34_port, S => q_2_0_34_port, Co => 
                           q_2_1_35_port);
   FA_C_1_0_35 : FA_551 port map( A => q_1_0_35_port, B => q_1_1_35_port, Ci =>
                           q_1_2_35_port, S => q_2_0_35_port, Co => 
                           q_2_1_36_port);
   FA_C_1_0_36 : FA_550 port map( A => q_1_0_36_port, B => q_1_1_36_port, Ci =>
                           q_1_2_36_port, S => q_2_0_36_port, Co => 
                           q_2_1_37_port);
   FA_C_1_0_37 : FA_549 port map( A => q_1_0_37_port, B => q_1_1_37_port, Ci =>
                           q_1_2_37_port, S => q_2_0_37_port, Co => 
                           q_2_1_38_port);
   FA_C_1_0_38 : FA_548 port map( A => q_1_0_38_port, B => q_1_1_38_port, Ci =>
                           q_1_2_38_port, S => q_2_0_38_port, Co => 
                           q_2_1_39_port);
   FA_C_1_0_39 : FA_547 port map( A => q_1_0_39_port, B => q_1_1_39_port, Ci =>
                           q_1_2_39_port, S => q_2_0_39_port, Co => 
                           q_2_1_40_port);
   FA_C_1_0_40 : FA_546 port map( A => q_1_0_40_port, B => q_1_1_40_port, Ci =>
                           q_1_2_40_port, S => q_2_0_40_port, Co => 
                           q_2_1_41_port);
   FA_C_1_0_41 : FA_545 port map( A => q_1_0_41_port, B => q_1_1_41_port, Ci =>
                           q_1_2_41_port, S => q_2_0_41_port, Co => 
                           q_2_1_42_port);
   FA_C_1_0_42 : FA_544 port map( A => q_1_0_42_port, B => q_1_1_42_port, Ci =>
                           q_0_2_42_port, S => q_2_0_42_port, Co => 
                           q_2_1_43_port);
   FA_C_1_0_43 : FA_543 port map( A => q_1_0_43_port, B => n91, Ci => 
                           q_0_1_43_port, S => q_2_0_43_port, Co => 
                           q_2_1_44_port);
   FA_C_1_0_44 : FA_542 port map( A => X_Logic1_port, B => q_0_1_44_port, Ci =>
                           q_0_2_44_port, S => q_2_0_44_port, Co => 
                           q_2_1_45_port);
   FA_C_1_0_45 : FA_541 port map( A => n90, B => q_0_1_45_port, Ci => 
                           q_0_2_45_port, S => q_2_0_45_port, Co => 
                           q_2_1_46_port);
   FA_C_1_0_46 : FA_540 port map( A => X_Logic1_port, B => q_0_1_46_port, Ci =>
                           q_0_2_46_port, S => q_2_0_46_port, Co => 
                           q_2_1_47_port);
   FA_C_1_0_47 : FA_539 port map( A => n89, B => q_0_1_47_port, Ci => 
                           q_0_2_47_port, S => q_2_0_47_port, Co => 
                           q_2_1_48_port);
   FA_C_1_0_48 : FA_538 port map( A => X_Logic1_port, B => q_0_1_48_port, Ci =>
                           q_0_2_48_port, S => q_2_0_48_port, Co => 
                           q_2_1_49_port);
   FA_C_1_0_49 : FA_537 port map( A => n88, B => q_0_1_49_port, Ci => 
                           q_0_2_49_port, S => q_2_0_49_port, Co => 
                           q_2_1_50_port);
   HA_L_1_0_50 : HA_30 port map( A => X_Logic1_port, B => q_0_1_50_port, S => 
                           q_2_0_50_port, C => q_2_0_51_port);
   HA_R_1_3_18 : HA_29 port map( A => q_0_3_18_port, B => q_0_4_18_port, S => 
                           q_2_2_18_port, C => q_2_3_19_port);
   HA_R_1_3_19 : HA_28 port map( A => q_0_3_19_port, B => q_0_4_19_port, S => 
                           q_2_2_19_port, C => q_2_3_20_port);
   FA_C_1_3_20 : FA_536 port map( A => q_0_3_20_port, B => q_0_4_20_port, Ci =>
                           q_0_5_20_port, S => q_2_2_20_port, Co => 
                           q_2_3_21_port);
   FA_C_1_3_21 : FA_535 port map( A => q_0_3_21_port, B => q_0_4_21_port, Ci =>
                           q_0_5_21_port, S => q_2_2_21_port, Co => 
                           q_2_3_22_port);
   FA_C_1_3_22 : FA_534 port map( A => q_0_3_22_port, B => q_0_4_22_port, Ci =>
                           q_0_5_22_port, S => q_2_2_22_port, Co => 
                           q_2_3_23_port);
   FA_C_1_3_23 : FA_533 port map( A => q_0_3_23_port, B => q_0_4_23_port, Ci =>
                           q_0_5_23_port, S => q_2_2_23_port, Co => 
                           q_2_3_24_port);
   FA_C_1_3_24 : FA_532 port map( A => q_0_4_24_port, B => q_0_5_24_port, Ci =>
                           q_0_6_24_port, S => q_2_2_24_port, Co => 
                           q_2_3_25_port);
   FA_C_1_3_25 : FA_531 port map( A => q_0_3_25_port, B => q_0_4_25_port, Ci =>
                           q_0_5_25_port, S => q_2_2_25_port, Co => 
                           q_2_3_26_port);
   FA_C_1_3_26 : FA_530 port map( A => q_0_5_26_port, B => q_0_6_26_port, Ci =>
                           q_0_7_26_port, S => q_2_2_26_port, Co => 
                           q_2_3_27_port);
   FA_C_1_3_27 : FA_529 port map( A => q_1_3_27_port, B => q_0_5_27_port, Ci =>
                           q_0_6_27_port, S => q_2_2_27_port, Co => 
                           q_2_3_28_port);
   FA_C_1_3_28 : FA_528 port map( A => q_1_3_28_port, B => q_1_4_28_port, Ci =>
                           q_0_8_28_port, S => q_2_2_28_port, Co => 
                           q_2_3_29_port);
   FA_C_1_3_29 : FA_527 port map( A => q_1_3_29_port, B => q_1_4_29_port, Ci =>
                           q_1_5_29_port, S => q_2_2_29_port, Co => 
                           q_2_3_30_port);
   FA_C_1_3_30 : FA_526 port map( A => q_1_3_30_port, B => q_1_4_30_port, Ci =>
                           q_1_5_30_port, S => q_2_2_30_port, Co => 
                           q_2_3_31_port);
   FA_C_1_3_31 : FA_525 port map( A => q_1_3_31_port, B => q_1_4_31_port, Ci =>
                           q_1_5_31_port, S => q_2_2_31_port, Co => 
                           q_2_3_32_port);
   FA_C_1_3_32 : FA_524 port map( A => q_1_3_32_port, B => q_1_4_32_port, Ci =>
                           q_1_5_32_port, S => q_2_2_32_port, Co => 
                           q_2_3_33_port);
   FA_C_1_3_33 : FA_523 port map( A => q_1_3_33_port, B => q_1_4_33_port, Ci =>
                           q_1_5_33_port, S => q_2_2_33_port, Co => 
                           q_2_3_34_port);
   FA_C_1_3_34 : FA_522 port map( A => q_1_3_34_port, B => q_1_4_34_port, Ci =>
                           q_1_5_34_port, S => q_2_2_34_port, Co => 
                           q_2_3_35_port);
   FA_C_1_3_35 : FA_521 port map( A => q_1_3_35_port, B => q_1_4_35_port, Ci =>
                           q_1_5_35_port, S => q_2_2_35_port, Co => 
                           q_2_3_36_port);
   FA_C_1_3_36 : FA_520 port map( A => q_1_3_36_port, B => q_1_4_36_port, Ci =>
                           q_1_5_36_port, S => q_2_2_36_port, Co => 
                           q_2_3_37_port);
   FA_C_1_3_37 : FA_519 port map( A => q_1_3_37_port, B => q_1_4_37_port, Ci =>
                           q_1_5_37_port, S => q_2_2_37_port, Co => 
                           q_2_3_38_port);
   FA_C_1_3_38 : FA_518 port map( A => q_1_3_38_port, B => q_1_4_38_port, Ci =>
                           q_1_5_38_port, S => q_2_2_38_port, Co => 
                           q_2_3_39_port);
   FA_C_1_3_39 : FA_517 port map( A => q_1_3_39_port, B => q_1_4_39_port, Ci =>
                           q_0_6_39_port, S => q_2_2_39_port, Co => 
                           q_2_3_40_port);
   FA_C_1_3_40 : FA_516 port map( A => q_1_3_40_port, B => q_0_5_40_port, Ci =>
                           q_0_6_40_port, S => q_2_2_40_port, Co => 
                           q_2_3_41_port);
   FA_C_1_3_41 : FA_515 port map( A => q_0_3_41_port, B => q_0_4_41_port, Ci =>
                           q_0_5_41_port, S => q_2_2_41_port, Co => 
                           q_2_3_42_port);
   FA_C_1_3_42 : FA_514 port map( A => q_0_3_42_port, B => q_0_4_42_port, Ci =>
                           q_0_5_42_port, S => q_2_2_42_port, Co => 
                           q_2_3_43_port);
   FA_C_1_3_43 : FA_513 port map( A => q_0_2_43_port, B => q_0_3_43_port, Ci =>
                           q_0_4_43_port, S => q_2_2_43_port, Co => 
                           q_2_3_44_port);
   FA_C_1_3_44 : FA_512 port map( A => q_0_3_44_port, B => q_0_4_44_port, Ci =>
                           q_0_5_44_port, S => q_2_2_44_port, Co => 
                           q_2_3_45_port);
   FA_C_1_3_45 : FA_511 port map( A => q_0_3_45_port, B => q_0_4_45_port, Ci =>
                           q_0_5_45_port, S => q_2_2_45_port, Co => 
                           q_2_3_46_port);
   FA_C_1_3_46 : FA_510 port map( A => q_0_3_46_port, B => q_0_4_46_port, Ci =>
                           q_0_5_46_port, S => q_2_2_46_port, Co => 
                           q_2_3_47_port);
   FA_C_1_3_47 : FA_509 port map( A => q_0_3_47_port, B => q_0_4_47_port, Ci =>
                           q_0_5_47_port, S => q_2_2_47_port, Co => 
                           q_2_3_48_port);
   HA_L_1_3_48 : HA_27 port map( A => q_0_3_48_port, B => q_0_4_48_port, S => 
                           q_2_2_48_port, C => q_2_2_49_port);
   HA_R_1_6_20 : HA_26 port map( A => q_0_6_20_port, B => q_0_7_20_port, S => 
                           q_2_4_20_port, C => q_2_5_21_port);
   HA_R_1_6_21 : HA_25 port map( A => q_0_6_21_port, B => q_0_7_21_port, S => 
                           q_2_4_21_port, C => q_2_5_22_port);
   FA_C_1_6_22 : FA_508 port map( A => q_0_6_22_port, B => q_0_7_22_port, Ci =>
                           q_0_8_22_port, S => q_2_4_22_port, Co => 
                           q_2_5_23_port);
   FA_C_1_6_23 : FA_507 port map( A => q_0_6_23_port, B => q_0_7_23_port, Ci =>
                           q_0_8_23_port, S => q_2_4_23_port, Co => 
                           q_2_5_24_port);
   FA_C_1_6_24 : FA_506 port map( A => q_0_7_24_port, B => q_0_8_24_port, Ci =>
                           q_0_9_24_port, S => q_2_4_24_port, Co => 
                           q_2_5_25_port);
   FA_C_1_6_25 : FA_505 port map( A => q_0_6_25_port, B => q_0_7_25_port, Ci =>
                           q_0_8_25_port, S => q_2_4_25_port, Co => 
                           q_2_5_26_port);
   FA_C_1_6_26 : FA_504 port map( A => q_0_8_26_port, B => q_0_9_26_port, Ci =>
                           q_0_10_26_port, S => q_2_4_26_port, Co => 
                           q_2_5_27_port);
   FA_C_1_6_27 : FA_503 port map( A => q_0_7_27_port, B => q_0_8_27_port, Ci =>
                           q_0_9_27_port, S => q_2_4_27_port, Co => 
                           q_2_5_28_port);
   FA_C_1_6_28 : FA_502 port map( A => q_0_9_28_port, B => q_0_10_28_port, Ci 
                           => q_0_11_28_port, S => q_2_4_28_port, Co => 
                           q_2_5_29_port);
   FA_C_1_6_29 : FA_501 port map( A => q_0_8_29_port, B => q_0_9_29_port, Ci =>
                           q_0_10_29_port, S => q_2_4_29_port, Co => 
                           q_2_5_30_port);
   FA_C_1_6_30 : FA_500 port map( A => q_1_6_30_port, B => q_0_11_30_port, Ci 
                           => q_0_12_30_port, S => q_2_4_30_port, Co => 
                           q_2_5_31_port);
   FA_C_1_6_31 : FA_499 port map( A => q_1_6_31_port, B => q_1_7_31_port, Ci =>
                           q_0_11_31_port, S => q_2_4_31_port, Co => 
                           q_2_5_32_port);
   FA_C_1_6_32 : FA_498 port map( A => q_1_6_32_port, B => q_1_7_32_port, Ci =>
                           q_0_12_32_port, S => q_2_4_32_port, Co => 
                           q_2_5_33_port);
   FA_C_1_6_33 : FA_497 port map( A => q_1_6_33_port, B => q_1_7_33_port, Ci =>
                           q_0_12_33_port, S => q_2_4_33_port, Co => 
                           q_2_5_34_port);
   FA_C_1_6_34 : FA_496 port map( A => q_1_6_34_port, B => q_1_7_34_port, Ci =>
                           q_0_12_34_port, S => q_2_4_34_port, Co => 
                           q_2_5_35_port);
   FA_C_1_6_35 : FA_495 port map( A => q_1_6_35_port, B => q_1_7_35_port, Ci =>
                           q_0_12_35_port, S => q_2_4_35_port, Co => 
                           q_2_5_36_port);
   FA_C_1_6_36 : FA_494 port map( A => q_1_6_36_port, B => q_1_7_36_port, Ci =>
                           q_0_11_36_port, S => q_2_4_36_port, Co => 
                           q_2_5_37_port);
   FA_C_1_6_37 : FA_493 port map( A => q_1_6_37_port, B => q_0_9_37_port, Ci =>
                           q_0_10_37_port, S => q_2_4_37_port, Co => 
                           q_2_5_38_port);
   FA_C_1_6_38 : FA_492 port map( A => q_0_8_38_port, B => q_0_9_38_port, Ci =>
                           q_0_10_38_port, S => q_2_4_38_port, Co => 
                           q_2_5_39_port);
   FA_C_1_6_39 : FA_491 port map( A => q_0_7_39_port, B => q_0_8_39_port, Ci =>
                           q_0_9_39_port, S => q_2_4_39_port, Co => 
                           q_2_5_40_port);
   FA_C_1_6_40 : FA_490 port map( A => q_0_7_40_port, B => q_0_8_40_port, Ci =>
                           q_0_9_40_port, S => q_2_4_40_port, Co => 
                           q_2_5_41_port);
   FA_C_1_6_41 : FA_489 port map( A => q_0_6_41_port, B => q_0_7_41_port, Ci =>
                           q_0_8_41_port, S => q_2_4_41_port, Co => 
                           q_2_5_42_port);
   FA_C_1_6_42 : FA_488 port map( A => q_0_6_42_port, B => q_0_7_42_port, Ci =>
                           q_0_8_42_port, S => q_2_4_42_port, Co => 
                           q_2_5_43_port);
   FA_C_1_6_43 : FA_487 port map( A => q_0_5_43_port, B => q_0_6_43_port, Ci =>
                           q_0_7_43_port, S => q_2_4_43_port, Co => 
                           q_2_5_44_port);
   FA_C_1_6_44 : FA_486 port map( A => q_0_6_44_port, B => q_0_7_44_port, Ci =>
                           q_0_8_44_port, S => q_2_4_44_port, Co => 
                           q_2_5_45_port);
   FA_C_1_6_45 : FA_485 port map( A => q_0_6_45_port, B => q_0_7_45_port, Ci =>
                           q_0_8_45_port, S => q_2_4_45_port, Co => 
                           q_2_5_46_port);
   HA_L_1_6_46 : HA_24 port map( A => q_0_6_46_port, B => q_0_7_46_port, S => 
                           q_2_4_46_port, C => q_2_4_47_port);
   HA_R_1_9_22 : HA_23 port map( A => q_0_9_22_port, B => q_0_10_22_port, S => 
                           q_2_6_22_port, C => q_2_7_23_port);
   HA_R_1_9_23 : HA_22 port map( A => q_0_9_23_port, B => q_0_10_23_port, S => 
                           q_2_6_23_port, C => q_2_7_24_port);
   FA_C_1_9_24 : FA_484 port map( A => q_0_10_24_port, B => q_0_11_24_port, Ci 
                           => q_0_12_24_port, S => q_2_6_24_port, Co => 
                           q_2_7_25_port);
   FA_C_1_9_25 : FA_483 port map( A => q_0_9_25_port, B => q_0_10_25_port, Ci 
                           => q_0_11_25_port, S => q_2_6_25_port, Co => 
                           q_2_7_26_port);
   FA_C_1_9_26 : FA_482 port map( A => q_0_11_26_port, B => q_0_12_26_port, Ci 
                           => q_0_13_26_port, S => q_2_6_26_port, Co => 
                           q_2_7_27_port);
   FA_C_1_9_27 : FA_481 port map( A => q_0_10_27_port, B => q_0_11_27_port, Ci 
                           => q_0_12_27_port, S => q_2_6_27_port, Co => 
                           q_2_7_28_port);
   FA_C_1_9_28 : FA_480 port map( A => q_0_12_28_port, B => q_0_13_28_port, Ci 
                           => q_0_14_28_port, S => q_2_6_28_port, Co => 
                           q_2_7_29_port);
   FA_C_1_9_29 : FA_479 port map( A => q_0_11_29_port, B => q_0_12_29_port, Ci 
                           => q_0_13_29_port, S => q_2_6_29_port, Co => 
                           q_2_7_30_port);
   FA_C_1_9_30 : FA_478 port map( A => q_0_13_30_port, B => q_0_14_30_port, Ci 
                           => q_0_15_30_port, S => q_2_6_30_port, Co => 
                           q_2_7_31_port);
   FA_C_1_9_31 : FA_477 port map( A => q_0_12_31_port, B => q_0_13_31_port, Ci 
                           => q_0_14_31_port, S => q_2_6_31_port, Co => 
                           q_2_7_32_port);
   FA_C_1_9_32 : FA_476 port map( A => q_0_13_32_port, B => q_0_14_32_port, Ci 
                           => q_0_15_32_port, S => q_2_6_32_port, Co => 
                           q_2_7_33_port);
   FA_C_1_9_33 : FA_475 port map( A => q_0_13_33_port, B => q_0_14_33_port, Ci 
                           => q_0_15_33_port, S => q_2_6_33_port, Co => 
                           q_2_7_34_port);
   FA_C_1_9_34 : FA_474 port map( A => q_0_13_34_port, B => q_0_14_34_port, Ci 
                           => q_0_15_34_port, S => q_2_6_34_port, Co => 
                           q_2_7_35_port);
   FA_C_1_9_35 : FA_473 port map( A => q_0_13_35_port, B => q_0_14_35_port, Ci 
                           => q_0_15_35_port, S => q_2_6_35_port, Co => 
                           q_2_7_36_port);
   FA_C_1_9_36 : FA_472 port map( A => q_0_12_36_port, B => q_0_13_36_port, Ci 
                           => q_0_14_36_port, S => q_2_6_36_port, Co => 
                           q_2_7_37_port);
   FA_C_1_9_37 : FA_471 port map( A => q_0_11_37_port, B => q_0_12_37_port, Ci 
                           => q_0_13_37_port, S => q_2_6_37_port, Co => 
                           q_2_7_38_port);
   FA_C_1_9_38 : FA_470 port map( A => q_0_11_38_port, B => q_0_12_38_port, Ci 
                           => q_0_13_38_port, S => q_2_6_38_port, Co => 
                           q_2_7_39_port);
   FA_C_1_9_39 : FA_469 port map( A => q_0_10_39_port, B => q_0_11_39_port, Ci 
                           => q_0_12_39_port, S => q_2_6_39_port, Co => 
                           q_2_7_40_port);
   FA_C_1_9_40 : FA_468 port map( A => q_0_10_40_port, B => q_0_11_40_port, Ci 
                           => q_0_12_40_port, S => q_2_6_40_port, Co => 
                           q_2_7_41_port);
   FA_C_1_9_41 : FA_467 port map( A => q_0_9_41_port, B => q_0_10_41_port, Ci 
                           => q_0_11_41_port, S => q_2_6_41_port, Co => 
                           q_2_7_42_port);
   FA_C_1_9_42 : FA_466 port map( A => q_0_9_42_port, B => q_0_10_42_port, Ci 
                           => q_0_11_42_port, S => q_2_6_42_port, Co => 
                           q_2_7_43_port);
   FA_C_1_9_43 : FA_465 port map( A => q_0_8_43_port, B => q_0_9_43_port, Ci =>
                           q_0_10_43_port, S => q_2_6_43_port, Co => 
                           q_2_7_44_port);
   HA_L_1_9_44 : HA_21 port map( A => q_0_9_44_port, B => q_0_10_44_port, S => 
                           q_2_6_44_port, C => q_2_6_45_port);
   HA_R_2_0_10 : HA_20 port map( A => q_0_0_10_port, B => q_0_1_10_port, S => 
                           q_3_0_10_port, C => q_3_1_11_port);
   HA_R_2_0_11 : HA_19 port map( A => q_0_0_11_port, B => q_0_1_11_port, S => 
                           q_3_0_11_port, C => q_3_1_12_port);
   FA_C_2_0_12 : FA_464 port map( A => q_0_0_12_port, B => q_0_1_12_port, Ci =>
                           q_0_2_12_port, S => q_3_0_12_port, Co => 
                           q_3_1_13_port);
   FA_C_2_0_13 : FA_463 port map( A => q_0_0_13_port, B => q_0_1_13_port, Ci =>
                           q_0_2_13_port, S => q_3_0_13_port, Co => 
                           q_3_1_14_port);
   FA_C_2_0_14 : FA_462 port map( A => q_0_0_14_port, B => q_0_1_14_port, Ci =>
                           q_0_2_14_port, S => q_3_0_14_port, Co => 
                           q_3_1_15_port);
   FA_C_2_0_15 : FA_461 port map( A => q_0_0_15_port, B => q_0_1_15_port, Ci =>
                           q_0_2_15_port, S => q_3_0_15_port, Co => 
                           q_3_1_16_port);
   FA_C_2_0_16 : FA_460 port map( A => q_2_0_16_port, B => q_0_2_16_port, Ci =>
                           q_0_3_16_port, S => q_3_0_16_port, Co => 
                           q_3_1_17_port);
   FA_C_2_0_17 : FA_459 port map( A => q_2_0_17_port, B => q_2_1_17_port, Ci =>
                           q_0_2_17_port, S => q_3_0_17_port, Co => 
                           q_3_1_18_port);
   FA_C_2_0_18 : FA_458 port map( A => q_2_0_18_port, B => q_2_1_18_port, Ci =>
                           q_2_2_18_port, S => q_3_0_18_port, Co => 
                           q_3_1_19_port);
   FA_C_2_0_19 : FA_457 port map( A => q_2_0_19_port, B => q_2_1_19_port, Ci =>
                           q_2_2_19_port, S => q_3_0_19_port, Co => 
                           q_3_1_20_port);
   FA_C_2_0_20 : FA_456 port map( A => q_2_0_20_port, B => q_2_1_20_port, Ci =>
                           q_2_2_20_port, S => q_3_0_20_port, Co => 
                           q_3_1_21_port);
   FA_C_2_0_21 : FA_455 port map( A => q_2_0_21_port, B => q_2_1_21_port, Ci =>
                           q_2_2_21_port, S => q_3_0_21_port, Co => 
                           q_3_1_22_port);
   FA_C_2_0_22 : FA_454 port map( A => q_2_0_22_port, B => q_2_1_22_port, Ci =>
                           q_2_2_22_port, S => q_3_0_22_port, Co => 
                           q_3_1_23_port);
   FA_C_2_0_23 : FA_453 port map( A => q_2_0_23_port, B => q_2_1_23_port, Ci =>
                           q_2_2_23_port, S => q_3_0_23_port, Co => 
                           q_3_1_24_port);
   FA_C_2_0_24 : FA_452 port map( A => q_2_0_24_port, B => q_2_1_24_port, Ci =>
                           q_2_2_24_port, S => q_3_0_24_port, Co => 
                           q_3_1_25_port);
   FA_C_2_0_25 : FA_451 port map( A => q_2_0_25_port, B => q_2_1_25_port, Ci =>
                           q_2_2_25_port, S => q_3_0_25_port, Co => 
                           q_3_1_26_port);
   FA_C_2_0_26 : FA_450 port map( A => q_2_0_26_port, B => q_2_1_26_port, Ci =>
                           q_2_2_26_port, S => q_3_0_26_port, Co => 
                           q_3_1_27_port);
   FA_C_2_0_27 : FA_449 port map( A => q_2_0_27_port, B => q_2_1_27_port, Ci =>
                           q_2_2_27_port, S => q_3_0_27_port, Co => 
                           q_3_1_28_port);
   FA_C_2_0_28 : FA_448 port map( A => q_2_0_28_port, B => q_2_1_28_port, Ci =>
                           q_2_2_28_port, S => q_3_0_28_port, Co => 
                           q_3_1_29_port);
   FA_C_2_0_29 : FA_447 port map( A => q_2_0_29_port, B => q_2_1_29_port, Ci =>
                           q_2_2_29_port, S => q_3_0_29_port, Co => 
                           q_3_1_30_port);
   FA_C_2_0_30 : FA_446 port map( A => q_2_0_30_port, B => q_2_1_30_port, Ci =>
                           q_2_2_30_port, S => q_3_0_30_port, Co => 
                           q_3_1_31_port);
   FA_C_2_0_31 : FA_445 port map( A => q_2_0_31_port, B => q_2_1_31_port, Ci =>
                           q_2_2_31_port, S => q_3_0_31_port, Co => 
                           q_3_1_32_port);
   FA_C_2_0_32 : FA_444 port map( A => q_2_0_32_port, B => q_2_1_32_port, Ci =>
                           q_2_2_32_port, S => q_3_0_32_port, Co => 
                           q_3_1_33_port);
   FA_C_2_0_33 : FA_443 port map( A => q_2_0_33_port, B => q_2_1_33_port, Ci =>
                           q_2_2_33_port, S => q_3_0_33_port, Co => 
                           q_3_1_34_port);
   FA_C_2_0_34 : FA_442 port map( A => q_2_0_34_port, B => q_2_1_34_port, Ci =>
                           q_2_2_34_port, S => q_3_0_34_port, Co => 
                           q_3_1_35_port);
   FA_C_2_0_35 : FA_441 port map( A => q_2_0_35_port, B => q_2_1_35_port, Ci =>
                           q_2_2_35_port, S => q_3_0_35_port, Co => 
                           q_3_1_36_port);
   FA_C_2_0_36 : FA_440 port map( A => q_2_0_36_port, B => q_2_1_36_port, Ci =>
                           q_2_2_36_port, S => q_3_0_36_port, Co => 
                           q_3_1_37_port);
   FA_C_2_0_37 : FA_439 port map( A => q_2_0_37_port, B => q_2_1_37_port, Ci =>
                           q_2_2_37_port, S => q_3_0_37_port, Co => 
                           q_3_1_38_port);
   FA_C_2_0_38 : FA_438 port map( A => q_2_0_38_port, B => q_2_1_38_port, Ci =>
                           q_2_2_38_port, S => q_3_0_38_port, Co => 
                           q_3_1_39_port);
   FA_C_2_0_39 : FA_437 port map( A => q_2_0_39_port, B => q_2_1_39_port, Ci =>
                           q_2_2_39_port, S => q_3_0_39_port, Co => 
                           q_3_1_40_port);
   FA_C_2_0_40 : FA_436 port map( A => q_2_0_40_port, B => q_2_1_40_port, Ci =>
                           q_2_2_40_port, S => q_3_0_40_port, Co => 
                           q_3_1_41_port);
   FA_C_2_0_41 : FA_435 port map( A => q_2_0_41_port, B => q_2_1_41_port, Ci =>
                           q_2_2_41_port, S => q_3_0_41_port, Co => 
                           q_3_1_42_port);
   FA_C_2_0_42 : FA_434 port map( A => q_2_0_42_port, B => q_2_1_42_port, Ci =>
                           q_2_2_42_port, S => q_3_0_42_port, Co => 
                           q_3_1_43_port);
   FA_C_2_0_43 : FA_433 port map( A => q_2_0_43_port, B => q_2_1_43_port, Ci =>
                           q_2_2_43_port, S => q_3_0_43_port, Co => 
                           q_3_1_44_port);
   FA_C_2_0_44 : FA_432 port map( A => q_2_0_44_port, B => q_2_1_44_port, Ci =>
                           q_2_2_44_port, S => q_3_0_44_port, Co => 
                           q_3_1_45_port);
   FA_C_2_0_45 : FA_431 port map( A => q_2_0_45_port, B => q_2_1_45_port, Ci =>
                           q_2_2_45_port, S => q_3_0_45_port, Co => 
                           q_3_1_46_port);
   FA_C_2_0_46 : FA_430 port map( A => q_2_0_46_port, B => q_2_1_46_port, Ci =>
                           q_2_2_46_port, S => q_3_0_46_port, Co => 
                           q_3_1_47_port);
   FA_C_2_0_47 : FA_429 port map( A => q_2_0_47_port, B => q_2_1_47_port, Ci =>
                           q_2_2_47_port, S => q_3_0_47_port, Co => 
                           q_3_1_48_port);
   FA_C_2_0_48 : FA_428 port map( A => q_2_0_48_port, B => q_2_1_48_port, Ci =>
                           q_2_2_48_port, S => q_3_0_48_port, Co => 
                           q_3_1_49_port);
   FA_C_2_0_49 : FA_427 port map( A => q_2_0_49_port, B => q_2_1_49_port, Ci =>
                           q_2_2_49_port, S => q_3_0_49_port, Co => 
                           q_3_1_50_port);
   FA_C_2_0_50 : FA_426 port map( A => q_2_0_50_port, B => q_2_1_50_port, Ci =>
                           q_0_2_50_port, S => q_3_0_50_port, Co => 
                           q_3_1_51_port);
   FA_C_2_0_51 : FA_425 port map( A => q_2_0_51_port, B => n87, Ci => 
                           q_0_1_51_port, S => q_3_0_51_port, Co => 
                           q_3_1_52_port);
   FA_C_2_0_52 : FA_424 port map( A => X_Logic1_port, B => q_0_1_52_port, Ci =>
                           q_0_2_52_port, S => q_3_0_52_port, Co => 
                           q_3_1_53_port);
   FA_C_2_0_53 : FA_423 port map( A => n86, B => q_0_1_53_port, Ci => 
                           q_0_2_53_port, S => q_3_0_53_port, Co => 
                           q_3_1_54_port);
   FA_C_2_0_54 : FA_422 port map( A => X_Logic1_port, B => q_0_1_54_port, Ci =>
                           q_0_2_54_port, S => q_3_0_54_port, Co => 
                           q_3_1_55_port);
   FA_C_2_0_55 : FA_421 port map( A => n85, B => q_0_1_55_port, Ci => 
                           q_0_2_55_port, S => q_3_0_55_port, Co => 
                           q_3_1_56_port);
   HA_L_2_0_56 : HA_18 port map( A => X_Logic1_port, B => q_0_1_56_port, S => 
                           q_3_0_56_port, C => q_3_0_57_port);
   HA_R_2_3_12 : HA_17 port map( A => q_0_3_12_port, B => q_0_4_12_port, S => 
                           q_3_2_12_port, C => q_3_3_13_port);
   HA_R_2_3_13 : HA_16 port map( A => q_0_3_13_port, B => q_0_4_13_port, S => 
                           q_3_2_13_port, C => q_3_3_14_port);
   FA_C_2_3_14 : FA_420 port map( A => q_0_3_14_port, B => q_0_4_14_port, Ci =>
                           q_0_5_14_port, S => q_3_2_14_port, Co => 
                           q_3_3_15_port);
   FA_C_2_3_15 : FA_419 port map( A => q_0_3_15_port, B => q_0_4_15_port, Ci =>
                           q_0_5_15_port, S => q_3_2_15_port, Co => 
                           q_3_3_16_port);
   FA_C_2_3_16 : FA_418 port map( A => q_0_4_16_port, B => q_0_5_16_port, Ci =>
                           q_0_6_16_port, S => q_3_2_16_port, Co => 
                           q_3_3_17_port);
   FA_C_2_3_17 : FA_417 port map( A => q_0_3_17_port, B => q_0_4_17_port, Ci =>
                           q_0_5_17_port, S => q_3_2_17_port, Co => 
                           q_3_3_18_port);
   FA_C_2_3_18 : FA_416 port map( A => q_0_5_18_port, B => q_0_6_18_port, Ci =>
                           q_0_7_18_port, S => q_3_2_18_port, Co => 
                           q_3_3_19_port);
   FA_C_2_3_19 : FA_415 port map( A => q_2_3_19_port, B => q_0_5_19_port, Ci =>
                           q_0_6_19_port, S => q_3_2_19_port, Co => 
                           q_3_3_20_port);
   FA_C_2_3_20 : FA_414 port map( A => q_2_3_20_port, B => q_2_4_20_port, Ci =>
                           q_0_8_20_port, S => q_3_2_20_port, Co => 
                           q_3_3_21_port);
   FA_C_2_3_21 : FA_413 port map( A => q_2_3_21_port, B => q_2_4_21_port, Ci =>
                           q_2_5_21_port, S => q_3_2_21_port, Co => 
                           q_3_3_22_port);
   FA_C_2_3_22 : FA_412 port map( A => q_2_3_22_port, B => q_2_4_22_port, Ci =>
                           q_2_5_22_port, S => q_3_2_22_port, Co => 
                           q_3_3_23_port);
   FA_C_2_3_23 : FA_411 port map( A => q_2_3_23_port, B => q_2_4_23_port, Ci =>
                           q_2_5_23_port, S => q_3_2_23_port, Co => 
                           q_3_3_24_port);
   FA_C_2_3_24 : FA_410 port map( A => q_2_3_24_port, B => q_2_4_24_port, Ci =>
                           q_2_5_24_port, S => q_3_2_24_port, Co => 
                           q_3_3_25_port);
   FA_C_2_3_25 : FA_409 port map( A => q_2_3_25_port, B => q_2_4_25_port, Ci =>
                           q_2_5_25_port, S => q_3_2_25_port, Co => 
                           q_3_3_26_port);
   FA_C_2_3_26 : FA_408 port map( A => q_2_3_26_port, B => q_2_4_26_port, Ci =>
                           q_2_5_26_port, S => q_3_2_26_port, Co => 
                           q_3_3_27_port);
   FA_C_2_3_27 : FA_407 port map( A => q_2_3_27_port, B => q_2_4_27_port, Ci =>
                           q_2_5_27_port, S => q_3_2_27_port, Co => 
                           q_3_3_28_port);
   FA_C_2_3_28 : FA_406 port map( A => q_2_3_28_port, B => q_2_4_28_port, Ci =>
                           q_2_5_28_port, S => q_3_2_28_port, Co => 
                           q_3_3_29_port);
   FA_C_2_3_29 : FA_405 port map( A => q_2_3_29_port, B => q_2_4_29_port, Ci =>
                           q_2_5_29_port, S => q_3_2_29_port, Co => 
                           q_3_3_30_port);
   FA_C_2_3_30 : FA_404 port map( A => q_2_3_30_port, B => q_2_4_30_port, Ci =>
                           q_2_5_30_port, S => q_3_2_30_port, Co => 
                           q_3_3_31_port);
   FA_C_2_3_31 : FA_403 port map( A => q_2_3_31_port, B => q_2_4_31_port, Ci =>
                           q_2_5_31_port, S => q_3_2_31_port, Co => 
                           q_3_3_32_port);
   FA_C_2_3_32 : FA_402 port map( A => q_2_3_32_port, B => q_2_4_32_port, Ci =>
                           q_2_5_32_port, S => q_3_2_32_port, Co => 
                           q_3_3_33_port);
   FA_C_2_3_33 : FA_401 port map( A => q_2_3_33_port, B => q_2_4_33_port, Ci =>
                           q_2_5_33_port, S => q_3_2_33_port, Co => 
                           q_3_3_34_port);
   FA_C_2_3_34 : FA_400 port map( A => q_2_3_34_port, B => q_2_4_34_port, Ci =>
                           q_2_5_34_port, S => q_3_2_34_port, Co => 
                           q_3_3_35_port);
   FA_C_2_3_35 : FA_399 port map( A => q_2_3_35_port, B => q_2_4_35_port, Ci =>
                           q_2_5_35_port, S => q_3_2_35_port, Co => 
                           q_3_3_36_port);
   FA_C_2_3_36 : FA_398 port map( A => q_2_3_36_port, B => q_2_4_36_port, Ci =>
                           q_2_5_36_port, S => q_3_2_36_port, Co => 
                           q_3_3_37_port);
   FA_C_2_3_37 : FA_397 port map( A => q_2_3_37_port, B => q_2_4_37_port, Ci =>
                           q_2_5_37_port, S => q_3_2_37_port, Co => 
                           q_3_3_38_port);
   FA_C_2_3_38 : FA_396 port map( A => q_2_3_38_port, B => q_2_4_38_port, Ci =>
                           q_2_5_38_port, S => q_3_2_38_port, Co => 
                           q_3_3_39_port);
   FA_C_2_3_39 : FA_395 port map( A => q_2_3_39_port, B => q_2_4_39_port, Ci =>
                           q_2_5_39_port, S => q_3_2_39_port, Co => 
                           q_3_3_40_port);
   FA_C_2_3_40 : FA_394 port map( A => q_2_3_40_port, B => q_2_4_40_port, Ci =>
                           q_2_5_40_port, S => q_3_2_40_port, Co => 
                           q_3_3_41_port);
   FA_C_2_3_41 : FA_393 port map( A => q_2_3_41_port, B => q_2_4_41_port, Ci =>
                           q_2_5_41_port, S => q_3_2_41_port, Co => 
                           q_3_3_42_port);
   FA_C_2_3_42 : FA_392 port map( A => q_2_3_42_port, B => q_2_4_42_port, Ci =>
                           q_2_5_42_port, S => q_3_2_42_port, Co => 
                           q_3_3_43_port);
   FA_C_2_3_43 : FA_391 port map( A => q_2_3_43_port, B => q_2_4_43_port, Ci =>
                           q_2_5_43_port, S => q_3_2_43_port, Co => 
                           q_3_3_44_port);
   FA_C_2_3_44 : FA_390 port map( A => q_2_3_44_port, B => q_2_4_44_port, Ci =>
                           q_2_5_44_port, S => q_3_2_44_port, Co => 
                           q_3_3_45_port);
   FA_C_2_3_45 : FA_389 port map( A => q_2_3_45_port, B => q_2_4_45_port, Ci =>
                           q_2_5_45_port, S => q_3_2_45_port, Co => 
                           q_3_3_46_port);
   FA_C_2_3_46 : FA_388 port map( A => q_2_3_46_port, B => q_2_4_46_port, Ci =>
                           q_2_5_46_port, S => q_3_2_46_port, Co => 
                           q_3_3_47_port);
   FA_C_2_3_47 : FA_387 port map( A => q_2_3_47_port, B => q_2_4_47_port, Ci =>
                           q_0_6_47_port, S => q_3_2_47_port, Co => 
                           q_3_3_48_port);
   FA_C_2_3_48 : FA_386 port map( A => q_2_3_48_port, B => q_0_5_48_port, Ci =>
                           q_0_6_48_port, S => q_3_2_48_port, Co => 
                           q_3_3_49_port);
   FA_C_2_3_49 : FA_385 port map( A => q_0_3_49_port, B => q_0_4_49_port, Ci =>
                           q_0_5_49_port, S => q_3_2_49_port, Co => 
                           q_3_3_50_port);
   FA_C_2_3_50 : FA_384 port map( A => q_0_3_50_port, B => q_0_4_50_port, Ci =>
                           q_0_5_50_port, S => q_3_2_50_port, Co => 
                           q_3_3_51_port);
   FA_C_2_3_51 : FA_383 port map( A => q_0_2_51_port, B => q_0_3_51_port, Ci =>
                           q_0_4_51_port, S => q_3_2_51_port, Co => 
                           q_3_3_52_port);
   FA_C_2_3_52 : FA_382 port map( A => q_0_3_52_port, B => q_0_4_52_port, Ci =>
                           q_0_5_52_port, S => q_3_2_52_port, Co => 
                           q_3_3_53_port);
   FA_C_2_3_53 : FA_381 port map( A => q_0_3_53_port, B => q_0_4_53_port, Ci =>
                           q_0_5_53_port, S => q_3_2_53_port, Co => 
                           q_3_3_54_port);
   HA_L_2_3_54 : HA_15 port map( A => q_0_3_54_port, B => q_0_4_54_port, S => 
                           q_3_2_54_port, C => q_3_2_55_port);
   HA_R_2_6_14 : HA_14 port map( A => q_0_6_14_port, B => q_0_7_14_port, S => 
                           q_3_4_14_port, C => q_3_5_15_port);
   HA_R_2_6_15 : HA_13 port map( A => q_0_6_15_port, B => q_0_7_15_port, S => 
                           q_3_4_15_port, C => q_3_5_16_port);
   FA_C_2_6_16 : FA_380 port map( A => q_0_7_16_port, B => q_0_8_16_port, Ci =>
                           n7, S => q_3_4_16_port, Co => q_3_5_17_port);
   FA_C_2_6_17 : FA_379 port map( A => q_0_6_17_port, B => q_0_7_17_port, Ci =>
                           q_0_8_17_port, S => q_3_4_17_port, Co => 
                           q_3_5_18_port);
   FA_C_2_6_18 : FA_378 port map( A => q_0_8_18_port, B => q_0_9_18_port, Ci =>
                           n9, S => q_3_4_18_port, Co => q_3_5_19_port);
   FA_C_2_6_19 : FA_377 port map( A => q_0_7_19_port, B => q_0_8_19_port, Ci =>
                           q_0_9_19_port, S => q_3_4_19_port, Co => 
                           q_3_5_20_port);
   FA_C_2_6_20 : FA_376 port map( A => q_0_9_20_port, B => q_0_10_20_port, Ci 
                           => n4, S => q_3_4_20_port, Co => q_3_5_21_port);
   FA_C_2_6_21 : FA_375 port map( A => q_0_8_21_port, B => q_0_9_21_port, Ci =>
                           q_0_10_21_port, S => q_3_4_21_port, Co => 
                           q_3_5_22_port);
   FA_C_2_6_22 : FA_374 port map( A => q_2_6_22_port, B => q_0_11_22_port, Ci 
                           => n6, S => q_3_4_22_port, Co => q_3_5_23_port);
   FA_C_2_6_23 : FA_373 port map( A => q_2_6_23_port, B => q_2_7_23_port, Ci =>
                           q_0_11_23_port, S => q_3_4_23_port, Co => 
                           q_3_5_24_port);
   FA_C_2_6_24 : FA_372 port map( A => q_2_6_24_port, B => q_2_7_24_port, Ci =>
                           B(25), S => q_3_4_24_port, Co => q_3_5_25_port);
   FA_C_2_6_25 : FA_371 port map( A => q_2_6_25_port, B => q_2_7_25_port, Ci =>
                           q_0_12_25_port, S => q_3_4_25_port, Co => 
                           q_3_5_26_port);
   FA_C_2_6_26 : FA_370 port map( A => q_2_6_26_port, B => q_2_7_26_port, Ci =>
                           B(27), S => q_3_4_26_port, Co => q_3_5_27_port);
   FA_C_2_6_27 : FA_369 port map( A => q_2_6_27_port, B => q_2_7_27_port, Ci =>
                           q_0_13_27_port, S => q_3_4_27_port, Co => 
                           q_3_5_28_port);
   FA_C_2_6_28 : FA_368 port map( A => q_2_6_28_port, B => q_2_7_28_port, Ci =>
                           B(29), S => q_3_4_28_port, Co => q_3_5_29_port);
   FA_C_2_6_29 : FA_367 port map( A => q_2_6_29_port, B => q_2_7_29_port, Ci =>
                           q_0_14_29_port, S => q_3_4_29_port, Co => 
                           q_3_5_30_port);
   FA_C_2_6_30 : FA_366 port map( A => q_2_6_30_port, B => q_2_7_30_port, Ci =>
                           B(31), S => q_3_4_30_port, Co => q_3_5_31_port);
   FA_C_2_6_31 : FA_365 port map( A => q_2_6_31_port, B => q_2_7_31_port, Ci =>
                           q_0_15_31_port, S => q_3_4_31_port, Co => 
                           q_3_5_32_port);
   FA_C_2_6_32 : FA_364 port map( A => q_2_6_32_port, B => q_2_7_32_port, Ci =>
                           q_0_16_32_port, S => q_3_4_32_port, Co => 
                           q_3_5_33_port);
   FA_C_2_6_33 : FA_363 port map( A => q_2_6_33_port, B => q_2_7_33_port, Ci =>
                           q_0_16_33_port, S => q_3_4_33_port, Co => 
                           q_3_5_34_port);
   FA_C_2_6_34 : FA_362 port map( A => q_2_6_34_port, B => q_2_7_34_port, Ci =>
                           q_0_16_34_port, S => q_3_4_34_port, Co => 
                           q_3_5_35_port);
   FA_C_2_6_35 : FA_361 port map( A => q_2_6_35_port, B => q_2_7_35_port, Ci =>
                           q_0_16_35_port, S => q_3_4_35_port, Co => 
                           q_3_5_36_port);
   FA_C_2_6_36 : FA_360 port map( A => q_2_6_36_port, B => q_2_7_36_port, Ci =>
                           q_0_15_36_port, S => q_3_4_36_port, Co => 
                           q_3_5_37_port);
   FA_C_2_6_37 : FA_359 port map( A => q_2_6_37_port, B => q_2_7_37_port, Ci =>
                           q_0_14_37_port, S => q_3_4_37_port, Co => 
                           q_3_5_38_port);
   FA_C_2_6_38 : FA_358 port map( A => q_2_6_38_port, B => q_2_7_38_port, Ci =>
                           q_0_14_38_port, S => q_3_4_38_port, Co => 
                           q_3_5_39_port);
   FA_C_2_6_39 : FA_357 port map( A => q_2_6_39_port, B => q_2_7_39_port, Ci =>
                           q_0_13_39_port, S => q_3_4_39_port, Co => 
                           q_3_5_40_port);
   FA_C_2_6_40 : FA_356 port map( A => q_2_6_40_port, B => q_2_7_40_port, Ci =>
                           q_0_13_40_port, S => q_3_4_40_port, Co => 
                           q_3_5_41_port);
   FA_C_2_6_41 : FA_355 port map( A => q_2_6_41_port, B => q_2_7_41_port, Ci =>
                           q_0_12_41_port, S => q_3_4_41_port, Co => 
                           q_3_5_42_port);
   FA_C_2_6_42 : FA_354 port map( A => q_2_6_42_port, B => q_2_7_42_port, Ci =>
                           q_0_12_42_port, S => q_3_4_42_port, Co => 
                           q_3_5_43_port);
   FA_C_2_6_43 : FA_353 port map( A => q_2_6_43_port, B => q_2_7_43_port, Ci =>
                           q_0_11_43_port, S => q_3_4_43_port, Co => 
                           q_3_5_44_port);
   FA_C_2_6_44 : FA_352 port map( A => q_2_6_44_port, B => q_2_7_44_port, Ci =>
                           q_0_11_44_port, S => q_3_4_44_port, Co => 
                           q_3_5_45_port);
   FA_C_2_6_45 : FA_351 port map( A => q_2_6_45_port, B => q_0_9_45_port, Ci =>
                           q_0_10_45_port, S => q_3_4_45_port, Co => 
                           q_3_5_46_port);
   FA_C_2_6_46 : FA_350 port map( A => q_0_8_46_port, B => q_0_9_46_port, Ci =>
                           q_0_10_46_port, S => q_3_4_46_port, Co => 
                           q_3_5_47_port);
   FA_C_2_6_47 : FA_349 port map( A => q_0_7_47_port, B => q_0_8_47_port, Ci =>
                           q_0_9_47_port, S => q_3_4_47_port, Co => 
                           q_3_5_48_port);
   FA_C_2_6_48 : FA_348 port map( A => q_0_7_48_port, B => q_0_8_48_port, Ci =>
                           q_0_9_48_port, S => q_3_4_48_port, Co => 
                           q_3_5_49_port);
   FA_C_2_6_49 : FA_347 port map( A => q_0_6_49_port, B => q_0_7_49_port, Ci =>
                           q_0_8_49_port, S => q_3_4_49_port, Co => 
                           q_3_5_50_port);
   FA_C_2_6_50 : FA_346 port map( A => q_0_6_50_port, B => q_0_7_50_port, Ci =>
                           q_0_8_50_port, S => q_3_4_50_port, Co => 
                           q_3_5_51_port);
   FA_C_2_6_51 : FA_345 port map( A => q_0_5_51_port, B => q_0_6_51_port, Ci =>
                           q_0_7_51_port, S => q_3_4_51_port, Co => 
                           q_3_5_52_port);
   HA_L_2_6_52 : HA_12 port map( A => q_0_6_52_port, B => q_0_7_52_port, S => 
                           q_3_4_52_port, C => q_3_4_53_port);
   HA_R_3_0_6 : HA_11 port map( A => q_0_0_6_port, B => q_0_1_6_port, S => 
                           q_4_0_6_port, C => q_4_1_7_port);
   HA_R_3_0_7 : HA_10 port map( A => q_0_0_7_port, B => q_0_1_7_port, S => 
                           q_4_0_7_port, C => q_4_1_8_port);
   FA_C_3_0_8 : FA_344 port map( A => q_0_0_8_port, B => q_0_1_8_port, Ci => 
                           q_0_2_8_port, S => q_4_0_8_port, Co => q_4_1_9_port)
                           ;
   FA_C_3_0_9 : FA_343 port map( A => q_0_0_9_port, B => q_0_1_9_port, Ci => 
                           q_0_2_9_port, S => q_4_0_9_port, Co => q_4_1_10_port
                           );
   FA_C_3_0_10 : FA_342 port map( A => q_3_0_10_port, B => q_0_2_10_port, Ci =>
                           q_0_3_10_port, S => q_4_0_10_port, Co => 
                           q_4_1_11_port);
   FA_C_3_0_11 : FA_341 port map( A => q_3_0_11_port, B => q_3_1_11_port, Ci =>
                           q_0_2_11_port, S => q_4_0_11_port, Co => 
                           q_4_1_12_port);
   FA_C_3_0_12 : FA_340 port map( A => q_3_0_12_port, B => q_3_1_12_port, Ci =>
                           q_3_2_12_port, S => q_4_0_12_port, Co => 
                           q_4_1_13_port);
   FA_C_3_0_13 : FA_339 port map( A => q_3_0_13_port, B => q_3_1_13_port, Ci =>
                           q_3_2_13_port, S => q_4_0_13_port, Co => 
                           q_4_1_14_port);
   FA_C_3_0_14 : FA_338 port map( A => q_3_0_14_port, B => q_3_1_14_port, Ci =>
                           q_3_2_14_port, S => q_4_0_14_port, Co => 
                           q_4_1_15_port);
   FA_C_3_0_15 : FA_337 port map( A => q_3_0_15_port, B => q_3_1_15_port, Ci =>
                           q_3_2_15_port, S => q_4_0_15_port, Co => 
                           q_4_1_16_port);
   FA_C_3_0_16 : FA_336 port map( A => q_3_0_16_port, B => q_3_1_16_port, Ci =>
                           q_3_2_16_port, S => q_4_0_16_port, Co => 
                           q_4_1_17_port);
   FA_C_3_0_17 : FA_335 port map( A => q_3_0_17_port, B => q_3_1_17_port, Ci =>
                           q_3_2_17_port, S => q_4_0_17_port, Co => 
                           q_4_1_18_port);
   FA_C_3_0_18 : FA_334 port map( A => q_3_0_18_port, B => q_3_1_18_port, Ci =>
                           q_3_2_18_port, S => q_4_0_18_port, Co => 
                           q_4_1_19_port);
   FA_C_3_0_19 : FA_333 port map( A => q_3_0_19_port, B => q_3_1_19_port, Ci =>
                           q_3_2_19_port, S => q_4_0_19_port, Co => 
                           q_4_1_20_port);
   FA_C_3_0_20 : FA_332 port map( A => q_3_0_20_port, B => q_3_1_20_port, Ci =>
                           q_3_2_20_port, S => q_4_0_20_port, Co => 
                           q_4_1_21_port);
   FA_C_3_0_21 : FA_331 port map( A => q_3_0_21_port, B => q_3_1_21_port, Ci =>
                           q_3_2_21_port, S => q_4_0_21_port, Co => 
                           q_4_1_22_port);
   FA_C_3_0_22 : FA_330 port map( A => q_3_0_22_port, B => q_3_1_22_port, Ci =>
                           q_3_2_22_port, S => q_4_0_22_port, Co => 
                           q_4_1_23_port);
   FA_C_3_0_23 : FA_329 port map( A => q_3_0_23_port, B => q_3_1_23_port, Ci =>
                           q_3_2_23_port, S => q_4_0_23_port, Co => 
                           q_4_1_24_port);
   FA_C_3_0_24 : FA_328 port map( A => q_3_0_24_port, B => q_3_1_24_port, Ci =>
                           q_3_2_24_port, S => q_4_0_24_port, Co => 
                           q_4_1_25_port);
   FA_C_3_0_25 : FA_327 port map( A => q_3_0_25_port, B => q_3_1_25_port, Ci =>
                           q_3_2_25_port, S => q_4_0_25_port, Co => 
                           q_4_1_26_port);
   FA_C_3_0_26 : FA_326 port map( A => q_3_0_26_port, B => q_3_1_26_port, Ci =>
                           q_3_2_26_port, S => q_4_0_26_port, Co => 
                           q_4_1_27_port);
   FA_C_3_0_27 : FA_325 port map( A => q_3_0_27_port, B => q_3_1_27_port, Ci =>
                           q_3_2_27_port, S => q_4_0_27_port, Co => 
                           q_4_1_28_port);
   FA_C_3_0_28 : FA_324 port map( A => q_3_0_28_port, B => q_3_1_28_port, Ci =>
                           q_3_2_28_port, S => q_4_0_28_port, Co => 
                           q_4_1_29_port);
   FA_C_3_0_29 : FA_323 port map( A => q_3_0_29_port, B => q_3_1_29_port, Ci =>
                           q_3_2_29_port, S => q_4_0_29_port, Co => 
                           q_4_1_30_port);
   FA_C_3_0_30 : FA_322 port map( A => q_3_0_30_port, B => q_3_1_30_port, Ci =>
                           q_3_2_30_port, S => q_4_0_30_port, Co => 
                           q_4_1_31_port);
   FA_C_3_0_31 : FA_321 port map( A => q_3_0_31_port, B => q_3_1_31_port, Ci =>
                           q_3_2_31_port, S => q_4_0_31_port, Co => 
                           q_4_1_32_port);
   FA_C_3_0_32 : FA_320 port map( A => q_3_0_32_port, B => q_3_1_32_port, Ci =>
                           q_3_2_32_port, S => q_4_0_32_port, Co => 
                           q_4_1_33_port);
   FA_C_3_0_33 : FA_319 port map( A => q_3_0_33_port, B => q_3_1_33_port, Ci =>
                           q_3_2_33_port, S => q_4_0_33_port, Co => 
                           q_4_1_34_port);
   FA_C_3_0_34 : FA_318 port map( A => q_3_0_34_port, B => q_3_1_34_port, Ci =>
                           q_3_2_34_port, S => q_4_0_34_port, Co => 
                           q_4_1_35_port);
   FA_C_3_0_35 : FA_317 port map( A => q_3_0_35_port, B => q_3_1_35_port, Ci =>
                           q_3_2_35_port, S => q_4_0_35_port, Co => 
                           q_4_1_36_port);
   FA_C_3_0_36 : FA_316 port map( A => q_3_0_36_port, B => q_3_1_36_port, Ci =>
                           q_3_2_36_port, S => q_4_0_36_port, Co => 
                           q_4_1_37_port);
   FA_C_3_0_37 : FA_315 port map( A => q_3_0_37_port, B => q_3_1_37_port, Ci =>
                           q_3_2_37_port, S => q_4_0_37_port, Co => 
                           q_4_1_38_port);
   FA_C_3_0_38 : FA_314 port map( A => q_3_0_38_port, B => q_3_1_38_port, Ci =>
                           q_3_2_38_port, S => q_4_0_38_port, Co => 
                           q_4_1_39_port);
   FA_C_3_0_39 : FA_313 port map( A => q_3_0_39_port, B => q_3_1_39_port, Ci =>
                           q_3_2_39_port, S => q_4_0_39_port, Co => 
                           q_4_1_40_port);
   FA_C_3_0_40 : FA_312 port map( A => q_3_0_40_port, B => q_3_1_40_port, Ci =>
                           q_3_2_40_port, S => q_4_0_40_port, Co => 
                           q_4_1_41_port);
   FA_C_3_0_41 : FA_311 port map( A => q_3_0_41_port, B => q_3_1_41_port, Ci =>
                           q_3_2_41_port, S => q_4_0_41_port, Co => 
                           q_4_1_42_port);
   FA_C_3_0_42 : FA_310 port map( A => q_3_0_42_port, B => q_3_1_42_port, Ci =>
                           q_3_2_42_port, S => q_4_0_42_port, Co => 
                           q_4_1_43_port);
   FA_C_3_0_43 : FA_309 port map( A => q_3_0_43_port, B => q_3_1_43_port, Ci =>
                           q_3_2_43_port, S => q_4_0_43_port, Co => 
                           q_4_1_44_port);
   FA_C_3_0_44 : FA_308 port map( A => q_3_0_44_port, B => q_3_1_44_port, Ci =>
                           q_3_2_44_port, S => q_4_0_44_port, Co => 
                           q_4_1_45_port);
   FA_C_3_0_45 : FA_307 port map( A => q_3_0_45_port, B => q_3_1_45_port, Ci =>
                           q_3_2_45_port, S => q_4_0_45_port, Co => 
                           q_4_1_46_port);
   FA_C_3_0_46 : FA_306 port map( A => q_3_0_46_port, B => q_3_1_46_port, Ci =>
                           q_3_2_46_port, S => q_4_0_46_port, Co => 
                           q_4_1_47_port);
   FA_C_3_0_47 : FA_305 port map( A => q_3_0_47_port, B => q_3_1_47_port, Ci =>
                           q_3_2_47_port, S => q_4_0_47_port, Co => 
                           q_4_1_48_port);
   FA_C_3_0_48 : FA_304 port map( A => q_3_0_48_port, B => q_3_1_48_port, Ci =>
                           q_3_2_48_port, S => q_4_0_48_port, Co => 
                           q_4_1_49_port);
   FA_C_3_0_49 : FA_303 port map( A => q_3_0_49_port, B => q_3_1_49_port, Ci =>
                           q_3_2_49_port, S => q_4_0_49_port, Co => 
                           q_4_1_50_port);
   FA_C_3_0_50 : FA_302 port map( A => q_3_0_50_port, B => q_3_1_50_port, Ci =>
                           q_3_2_50_port, S => q_4_0_50_port, Co => 
                           q_4_1_51_port);
   FA_C_3_0_51 : FA_301 port map( A => q_3_0_51_port, B => q_3_1_51_port, Ci =>
                           q_3_2_51_port, S => q_4_0_51_port, Co => 
                           q_4_1_52_port);
   FA_C_3_0_52 : FA_300 port map( A => q_3_0_52_port, B => q_3_1_52_port, Ci =>
                           q_3_2_52_port, S => q_4_0_52_port, Co => 
                           q_4_1_53_port);
   FA_C_3_0_53 : FA_299 port map( A => q_3_0_53_port, B => q_3_1_53_port, Ci =>
                           q_3_2_53_port, S => q_4_0_53_port, Co => 
                           q_4_1_54_port);
   FA_C_3_0_54 : FA_298 port map( A => q_3_0_54_port, B => q_3_1_54_port, Ci =>
                           q_3_2_54_port, S => q_4_0_54_port, Co => 
                           q_4_1_55_port);
   FA_C_3_0_55 : FA_297 port map( A => q_3_0_55_port, B => q_3_1_55_port, Ci =>
                           q_3_2_55_port, S => q_4_0_55_port, Co => 
                           q_4_1_56_port);
   FA_C_3_0_56 : FA_296 port map( A => q_3_0_56_port, B => q_3_1_56_port, Ci =>
                           q_0_2_56_port, S => q_4_0_56_port, Co => 
                           q_4_1_57_port);
   FA_C_3_0_57 : FA_295 port map( A => q_3_0_57_port, B => n84, Ci => 
                           q_0_1_57_port, S => q_4_0_57_port, Co => 
                           q_4_1_58_port);
   FA_C_3_0_58 : FA_294 port map( A => X_Logic1_port, B => q_0_1_58_port, Ci =>
                           q_0_2_58_port, S => q_4_0_58_port, Co => 
                           q_4_1_59_port);
   FA_C_3_0_59 : FA_293 port map( A => n83, B => q_0_1_59_port, Ci => 
                           q_0_2_59_port, S => q_4_0_59_port, Co => 
                           q_4_1_60_port);
   HA_L_3_0_60 : HA_9 port map( A => X_Logic1_port, B => q_0_1_60_port, S => 
                           q_4_0_60_port, C => q_4_0_61_port);
   HA_R_3_3_8 : HA_8 port map( A => q_0_3_8_port, B => q_0_4_8_port, S => 
                           q_4_2_8_port, C => q_5_2_9_port);
   HA_R_3_3_9 : HA_7 port map( A => q_0_3_9_port, B => q_0_4_9_port, S => 
                           q_4_2_9_port, C => q_5_2_10_port);
   FA_C_3_3_10 : FA_292 port map( A => q_0_4_10_port, B => q_0_5_10_port, Ci =>
                           n5, S => q_4_2_10_port, Co => q_5_2_11_port);
   FA_C_3_3_11 : FA_291 port map( A => q_0_3_11_port, B => q_0_4_11_port, Ci =>
                           q_0_5_11_port, S => q_4_2_11_port, Co => 
                           q_5_2_12_port);
   FA_C_3_3_12 : FA_290 port map( A => q_0_5_12_port, B => q_0_6_12_port, Ci =>
                           n1, S => q_4_2_12_port, Co => q_5_2_13_port);
   FA_C_3_3_13 : FA_289 port map( A => q_3_3_13_port, B => q_0_5_13_port, Ci =>
                           q_0_6_13_port, S => q_4_2_13_port, Co => 
                           q_5_2_14_port);
   FA_C_3_3_14 : FA_288 port map( A => q_3_3_14_port, B => q_3_4_14_port, Ci =>
                           n13, S => q_4_2_14_port, Co => q_5_2_15_port);
   FA_C_3_3_15 : FA_287 port map( A => q_3_3_15_port, B => q_3_4_15_port, Ci =>
                           q_3_5_15_port, S => q_4_2_15_port, Co => 
                           q_5_2_16_port);
   FA_C_3_3_16 : FA_286 port map( A => q_3_3_16_port, B => q_3_4_16_port, Ci =>
                           q_3_5_16_port, S => q_4_2_16_port, Co => 
                           q_5_2_17_port);
   FA_C_3_3_17 : FA_285 port map( A => q_3_3_17_port, B => q_3_4_17_port, Ci =>
                           q_3_5_17_port, S => q_4_2_17_port, Co => 
                           q_5_2_18_port);
   FA_C_3_3_18 : FA_284 port map( A => q_3_3_18_port, B => q_3_4_18_port, Ci =>
                           q_3_5_18_port, S => q_4_2_18_port, Co => 
                           q_5_2_19_port);
   FA_C_3_3_19 : FA_283 port map( A => q_3_3_19_port, B => q_3_4_19_port, Ci =>
                           q_3_5_19_port, S => q_4_2_19_port, Co => 
                           q_5_2_20_port);
   FA_C_3_3_20 : FA_282 port map( A => q_3_3_20_port, B => q_3_4_20_port, Ci =>
                           q_3_5_20_port, S => q_4_2_20_port, Co => 
                           q_5_2_21_port);
   FA_C_3_3_21 : FA_281 port map( A => q_3_3_21_port, B => q_3_4_21_port, Ci =>
                           q_3_5_21_port, S => q_4_2_21_port, Co => 
                           q_5_2_22_port);
   FA_C_3_3_22 : FA_280 port map( A => q_3_3_22_port, B => q_3_4_22_port, Ci =>
                           q_3_5_22_port, S => q_4_2_22_port, Co => 
                           q_5_2_23_port);
   FA_C_3_3_23 : FA_279 port map( A => q_3_3_23_port, B => q_3_4_23_port, Ci =>
                           q_3_5_23_port, S => q_4_2_23_port, Co => 
                           q_5_2_24_port);
   FA_C_3_3_24 : FA_278 port map( A => q_3_3_24_port, B => q_3_4_24_port, Ci =>
                           q_3_5_24_port, S => q_4_2_24_port, Co => 
                           q_5_2_25_port);
   FA_C_3_3_25 : FA_277 port map( A => q_3_3_25_port, B => q_3_4_25_port, Ci =>
                           q_3_5_25_port, S => q_4_2_25_port, Co => 
                           q_5_2_26_port);
   FA_C_3_3_26 : FA_276 port map( A => q_3_3_26_port, B => q_3_4_26_port, Ci =>
                           q_3_5_26_port, S => q_4_2_26_port, Co => 
                           q_5_2_27_port);
   FA_C_3_3_27 : FA_275 port map( A => q_3_3_27_port, B => q_3_4_27_port, Ci =>
                           q_3_5_27_port, S => q_4_2_27_port, Co => 
                           q_5_2_28_port);
   FA_C_3_3_28 : FA_274 port map( A => q_3_3_28_port, B => q_3_4_28_port, Ci =>
                           q_3_5_28_port, S => q_4_2_28_port, Co => 
                           q_5_2_29_port);
   FA_C_3_3_29 : FA_273 port map( A => q_3_3_29_port, B => q_3_4_29_port, Ci =>
                           q_3_5_29_port, S => q_4_2_29_port, Co => 
                           q_5_2_30_port);
   FA_C_3_3_30 : FA_272 port map( A => q_3_3_30_port, B => q_3_4_30_port, Ci =>
                           q_3_5_30_port, S => q_4_2_30_port, Co => 
                           q_5_2_31_port);
   FA_C_3_3_31 : FA_271 port map( A => q_3_3_31_port, B => q_3_4_31_port, Ci =>
                           q_3_5_31_port, S => q_4_2_31_port, Co => 
                           q_5_2_32_port);
   FA_C_3_3_32 : FA_270 port map( A => q_3_3_32_port, B => q_3_4_32_port, Ci =>
                           q_3_5_32_port, S => q_4_2_32_port, Co => 
                           q_5_2_33_port);
   FA_C_3_3_33 : FA_269 port map( A => q_3_3_33_port, B => q_3_4_33_port, Ci =>
                           q_3_5_33_port, S => q_4_2_33_port, Co => 
                           q_5_2_34_port);
   FA_C_3_3_34 : FA_268 port map( A => q_3_3_34_port, B => q_3_4_34_port, Ci =>
                           q_3_5_34_port, S => q_4_2_34_port, Co => 
                           q_5_2_35_port);
   FA_C_3_3_35 : FA_267 port map( A => q_3_3_35_port, B => q_3_4_35_port, Ci =>
                           q_3_5_35_port, S => q_4_2_35_port, Co => 
                           q_5_2_36_port);
   FA_C_3_3_36 : FA_266 port map( A => q_3_3_36_port, B => q_3_4_36_port, Ci =>
                           q_3_5_36_port, S => q_4_2_36_port, Co => 
                           q_5_2_37_port);
   FA_C_3_3_37 : FA_265 port map( A => q_3_3_37_port, B => q_3_4_37_port, Ci =>
                           q_3_5_37_port, S => q_4_2_37_port, Co => 
                           q_5_2_38_port);
   FA_C_3_3_38 : FA_264 port map( A => q_3_3_38_port, B => q_3_4_38_port, Ci =>
                           q_3_5_38_port, S => q_4_2_38_port, Co => 
                           q_5_2_39_port);
   FA_C_3_3_39 : FA_263 port map( A => q_3_3_39_port, B => q_3_4_39_port, Ci =>
                           q_3_5_39_port, S => q_4_2_39_port, Co => 
                           q_5_2_40_port);
   FA_C_3_3_40 : FA_262 port map( A => q_3_3_40_port, B => q_3_4_40_port, Ci =>
                           q_3_5_40_port, S => q_4_2_40_port, Co => 
                           q_5_2_41_port);
   FA_C_3_3_41 : FA_261 port map( A => q_3_3_41_port, B => q_3_4_41_port, Ci =>
                           q_3_5_41_port, S => q_4_2_41_port, Co => 
                           q_5_2_42_port);
   FA_C_3_3_42 : FA_260 port map( A => q_3_3_42_port, B => q_3_4_42_port, Ci =>
                           q_3_5_42_port, S => q_4_2_42_port, Co => 
                           q_5_2_43_port);
   FA_C_3_3_43 : FA_259 port map( A => q_3_3_43_port, B => q_3_4_43_port, Ci =>
                           q_3_5_43_port, S => q_4_2_43_port, Co => 
                           q_5_2_44_port);
   FA_C_3_3_44 : FA_258 port map( A => q_3_3_44_port, B => q_3_4_44_port, Ci =>
                           q_3_5_44_port, S => q_4_2_44_port, Co => 
                           q_5_2_45_port);
   FA_C_3_3_45 : FA_257 port map( A => q_3_3_45_port, B => q_3_4_45_port, Ci =>
                           q_3_5_45_port, S => q_4_2_45_port, Co => 
                           q_5_2_46_port);
   FA_C_3_3_46 : FA_256 port map( A => q_3_3_46_port, B => q_3_4_46_port, Ci =>
                           q_3_5_46_port, S => q_4_2_46_port, Co => 
                           q_5_2_47_port);
   FA_C_3_3_47 : FA_255 port map( A => q_3_3_47_port, B => q_3_4_47_port, Ci =>
                           q_3_5_47_port, S => q_4_2_47_port, Co => 
                           q_5_2_48_port);
   FA_C_3_3_48 : FA_254 port map( A => q_3_3_48_port, B => q_3_4_48_port, Ci =>
                           q_3_5_48_port, S => q_4_2_48_port, Co => 
                           q_5_2_49_port);
   FA_C_3_3_49 : FA_253 port map( A => q_3_3_49_port, B => q_3_4_49_port, Ci =>
                           q_3_5_49_port, S => q_4_2_49_port, Co => 
                           q_5_2_50_port);
   FA_C_3_3_50 : FA_252 port map( A => q_3_3_50_port, B => q_3_4_50_port, Ci =>
                           q_3_5_50_port, S => q_4_2_50_port, Co => 
                           q_5_2_51_port);
   FA_C_3_3_51 : FA_251 port map( A => q_3_3_51_port, B => q_3_4_51_port, Ci =>
                           q_3_5_51_port, S => q_4_2_51_port, Co => 
                           q_5_2_52_port);
   FA_C_3_3_52 : FA_250 port map( A => q_3_3_52_port, B => q_3_4_52_port, Ci =>
                           q_3_5_52_port, S => q_4_2_52_port, Co => 
                           q_5_2_53_port);
   FA_C_3_3_53 : FA_249 port map( A => q_3_3_53_port, B => q_3_4_53_port, Ci =>
                           q_0_6_53_port, S => q_4_2_53_port, Co => 
                           q_5_2_54_port);
   FA_C_3_3_54 : FA_248 port map( A => q_3_3_54_port, B => q_0_5_54_port, Ci =>
                           q_0_6_54_port, S => q_4_2_54_port, Co => 
                           q_5_2_55_port);
   FA_C_3_3_55 : FA_247 port map( A => q_0_3_55_port, B => q_0_4_55_port, Ci =>
                           q_0_5_55_port, S => q_4_2_55_port, Co => 
                           q_5_2_56_port);
   FA_C_3_3_56 : FA_246 port map( A => q_0_3_56_port, B => q_0_4_56_port, Ci =>
                           q_0_5_56_port, S => q_4_2_56_port, Co => 
                           q_5_2_57_port);
   FA_C_3_3_57 : FA_245 port map( A => q_0_2_57_port, B => q_0_3_57_port, Ci =>
                           q_0_4_57_port, S => q_4_2_57_port, Co => 
                           q_5_2_58_port);
   HA_L_3_3_58 : HA_6 port map( A => q_0_3_58_port, B => q_0_4_58_port, S => 
                           q_4_2_58_port, C => q_4_2_59_port);
   HA_R_4_0_4 : HA_5 port map( A => q_0_0_4_port, B => q_0_1_4_port, S => 
                           q_5_0_4_port, C => q_5_1_5_port);
   HA_R_4_0_5 : HA_4 port map( A => q_0_0_5_port, B => q_0_1_5_port, S => 
                           q_5_0_5_port, C => q_5_1_6_port);
   FA_C_4_0_6 : FA_244 port map( A => q_4_0_6_port, B => q_0_2_6_port, Ci => 
                           q_0_3_6_port, S => q_5_0_6_port, Co => q_5_1_7_port)
                           ;
   FA_C_4_0_7 : FA_243 port map( A => q_4_0_7_port, B => q_4_1_7_port, Ci => 
                           q_0_2_7_port, S => q_5_0_7_port, Co => q_5_1_8_port)
                           ;
   FA_C_4_0_8 : FA_242 port map( A => q_4_0_8_port, B => q_4_1_8_port, Ci => 
                           q_4_2_8_port, S => q_5_0_8_port, Co => q_5_1_9_port)
                           ;
   FA_C_4_0_9 : FA_241 port map( A => q_4_0_9_port, B => q_4_1_9_port, Ci => 
                           q_4_2_9_port, S => q_5_0_9_port, Co => q_5_1_10_port
                           );
   FA_C_4_0_10 : FA_240 port map( A => q_4_0_10_port, B => q_4_1_10_port, Ci =>
                           q_4_2_10_port, S => q_5_0_10_port, Co => 
                           q_5_1_11_port);
   FA_C_4_0_11 : FA_239 port map( A => q_4_0_11_port, B => q_4_1_11_port, Ci =>
                           q_4_2_11_port, S => q_5_0_11_port, Co => 
                           q_5_1_12_port);
   FA_C_4_0_12 : FA_238 port map( A => q_4_0_12_port, B => q_4_1_12_port, Ci =>
                           q_4_2_12_port, S => q_5_0_12_port, Co => 
                           q_5_1_13_port);
   FA_C_4_0_13 : FA_237 port map( A => q_4_0_13_port, B => q_4_1_13_port, Ci =>
                           q_4_2_13_port, S => q_5_0_13_port, Co => 
                           q_5_1_14_port);
   FA_C_4_0_14 : FA_236 port map( A => q_4_0_14_port, B => q_4_1_14_port, Ci =>
                           q_4_2_14_port, S => q_5_0_14_port, Co => 
                           q_5_1_15_port);
   FA_C_4_0_15 : FA_235 port map( A => q_4_0_15_port, B => q_4_1_15_port, Ci =>
                           q_4_2_15_port, S => q_5_0_15_port, Co => 
                           q_5_1_16_port);
   FA_C_4_0_16 : FA_234 port map( A => q_4_0_16_port, B => q_4_1_16_port, Ci =>
                           q_4_2_16_port, S => q_5_0_16_port, Co => 
                           q_5_1_17_port);
   FA_C_4_0_17 : FA_233 port map( A => q_4_0_17_port, B => q_4_1_17_port, Ci =>
                           q_4_2_17_port, S => q_5_0_17_port, Co => 
                           q_5_1_18_port);
   FA_C_4_0_18 : FA_232 port map( A => q_4_0_18_port, B => q_4_1_18_port, Ci =>
                           q_4_2_18_port, S => q_5_0_18_port, Co => 
                           q_5_1_19_port);
   FA_C_4_0_19 : FA_231 port map( A => q_4_0_19_port, B => q_4_1_19_port, Ci =>
                           q_4_2_19_port, S => q_5_0_19_port, Co => 
                           q_5_1_20_port);
   FA_C_4_0_20 : FA_230 port map( A => q_4_0_20_port, B => q_4_1_20_port, Ci =>
                           q_4_2_20_port, S => q_5_0_20_port, Co => 
                           q_5_1_21_port);
   FA_C_4_0_21 : FA_229 port map( A => q_4_0_21_port, B => q_4_1_21_port, Ci =>
                           q_4_2_21_port, S => q_5_0_21_port, Co => 
                           q_5_1_22_port);
   FA_C_4_0_22 : FA_228 port map( A => q_4_0_22_port, B => q_4_1_22_port, Ci =>
                           q_4_2_22_port, S => q_5_0_22_port, Co => 
                           q_5_1_23_port);
   FA_C_4_0_23 : FA_227 port map( A => q_4_0_23_port, B => q_4_1_23_port, Ci =>
                           q_4_2_23_port, S => q_5_0_23_port, Co => 
                           q_5_1_24_port);
   FA_C_4_0_24 : FA_226 port map( A => q_4_0_24_port, B => q_4_1_24_port, Ci =>
                           q_4_2_24_port, S => q_5_0_24_port, Co => 
                           q_5_1_25_port);
   FA_C_4_0_25 : FA_225 port map( A => q_4_0_25_port, B => q_4_1_25_port, Ci =>
                           q_4_2_25_port, S => q_5_0_25_port, Co => 
                           q_5_1_26_port);
   FA_C_4_0_26 : FA_224 port map( A => q_4_0_26_port, B => q_4_1_26_port, Ci =>
                           q_4_2_26_port, S => q_5_0_26_port, Co => 
                           q_5_1_27_port);
   FA_C_4_0_27 : FA_223 port map( A => q_4_0_27_port, B => q_4_1_27_port, Ci =>
                           q_4_2_27_port, S => q_5_0_27_port, Co => 
                           q_5_1_28_port);
   FA_C_4_0_28 : FA_222 port map( A => q_4_0_28_port, B => q_4_1_28_port, Ci =>
                           q_4_2_28_port, S => q_5_0_28_port, Co => 
                           q_5_1_29_port);
   FA_C_4_0_29 : FA_221 port map( A => q_4_0_29_port, B => q_4_1_29_port, Ci =>
                           q_4_2_29_port, S => q_5_0_29_port, Co => 
                           q_5_1_30_port);
   FA_C_4_0_30 : FA_220 port map( A => q_4_0_30_port, B => q_4_1_30_port, Ci =>
                           q_4_2_30_port, S => q_5_0_30_port, Co => 
                           q_5_1_31_port);
   FA_C_4_0_31 : FA_219 port map( A => q_4_0_31_port, B => q_4_1_31_port, Ci =>
                           q_4_2_31_port, S => q_5_0_31_port, Co => 
                           q_5_1_32_port);
   FA_C_4_0_32 : FA_218 port map( A => q_4_0_32_port, B => q_4_1_32_port, Ci =>
                           q_4_2_32_port, S => q_5_0_32_port, Co => 
                           q_5_1_33_port);
   FA_C_4_0_33 : FA_217 port map( A => q_4_0_33_port, B => q_4_1_33_port, Ci =>
                           q_4_2_33_port, S => q_5_0_33_port, Co => 
                           q_5_1_34_port);
   FA_C_4_0_34 : FA_216 port map( A => q_4_0_34_port, B => q_4_1_34_port, Ci =>
                           q_4_2_34_port, S => q_5_0_34_port, Co => 
                           q_5_1_35_port);
   FA_C_4_0_35 : FA_215 port map( A => q_4_0_35_port, B => q_4_1_35_port, Ci =>
                           q_4_2_35_port, S => q_5_0_35_port, Co => 
                           q_5_1_36_port);
   FA_C_4_0_36 : FA_214 port map( A => q_4_0_36_port, B => q_4_1_36_port, Ci =>
                           q_4_2_36_port, S => q_5_0_36_port, Co => 
                           q_5_1_37_port);
   FA_C_4_0_37 : FA_213 port map( A => q_4_0_37_port, B => q_4_1_37_port, Ci =>
                           q_4_2_37_port, S => q_5_0_37_port, Co => 
                           q_5_1_38_port);
   FA_C_4_0_38 : FA_212 port map( A => q_4_0_38_port, B => q_4_1_38_port, Ci =>
                           q_4_2_38_port, S => q_5_0_38_port, Co => 
                           q_5_1_39_port);
   FA_C_4_0_39 : FA_211 port map( A => q_4_0_39_port, B => q_4_1_39_port, Ci =>
                           q_4_2_39_port, S => q_5_0_39_port, Co => 
                           q_5_1_40_port);
   FA_C_4_0_40 : FA_210 port map( A => q_4_0_40_port, B => q_4_1_40_port, Ci =>
                           q_4_2_40_port, S => q_5_0_40_port, Co => 
                           q_5_1_41_port);
   FA_C_4_0_41 : FA_209 port map( A => q_4_0_41_port, B => q_4_1_41_port, Ci =>
                           q_4_2_41_port, S => q_5_0_41_port, Co => 
                           q_5_1_42_port);
   FA_C_4_0_42 : FA_208 port map( A => q_4_0_42_port, B => q_4_1_42_port, Ci =>
                           q_4_2_42_port, S => q_5_0_42_port, Co => 
                           q_5_1_43_port);
   FA_C_4_0_43 : FA_207 port map( A => q_4_0_43_port, B => q_4_1_43_port, Ci =>
                           q_4_2_43_port, S => q_5_0_43_port, Co => 
                           q_5_1_44_port);
   FA_C_4_0_44 : FA_206 port map( A => q_4_0_44_port, B => q_4_1_44_port, Ci =>
                           q_4_2_44_port, S => q_5_0_44_port, Co => 
                           q_5_1_45_port);
   FA_C_4_0_45 : FA_205 port map( A => q_4_0_45_port, B => q_4_1_45_port, Ci =>
                           q_4_2_45_port, S => q_5_0_45_port, Co => 
                           q_5_1_46_port);
   FA_C_4_0_46 : FA_204 port map( A => q_4_0_46_port, B => q_4_1_46_port, Ci =>
                           q_4_2_46_port, S => q_5_0_46_port, Co => 
                           q_5_1_47_port);
   FA_C_4_0_47 : FA_203 port map( A => q_4_0_47_port, B => q_4_1_47_port, Ci =>
                           q_4_2_47_port, S => q_5_0_47_port, Co => 
                           q_5_1_48_port);
   FA_C_4_0_48 : FA_202 port map( A => q_4_0_48_port, B => q_4_1_48_port, Ci =>
                           q_4_2_48_port, S => q_5_0_48_port, Co => 
                           q_5_1_49_port);
   FA_C_4_0_49 : FA_201 port map( A => q_4_0_49_port, B => q_4_1_49_port, Ci =>
                           q_4_2_49_port, S => q_5_0_49_port, Co => 
                           q_5_1_50_port);
   FA_C_4_0_50 : FA_200 port map( A => q_4_0_50_port, B => q_4_1_50_port, Ci =>
                           q_4_2_50_port, S => q_5_0_50_port, Co => 
                           q_5_1_51_port);
   FA_C_4_0_51 : FA_199 port map( A => q_4_0_51_port, B => q_4_1_51_port, Ci =>
                           q_4_2_51_port, S => q_5_0_51_port, Co => 
                           q_5_1_52_port);
   FA_C_4_0_52 : FA_198 port map( A => q_4_0_52_port, B => q_4_1_52_port, Ci =>
                           q_4_2_52_port, S => q_5_0_52_port, Co => 
                           q_5_1_53_port);
   FA_C_4_0_53 : FA_197 port map( A => q_4_0_53_port, B => q_4_1_53_port, Ci =>
                           q_4_2_53_port, S => q_5_0_53_port, Co => 
                           q_5_1_54_port);
   FA_C_4_0_54 : FA_196 port map( A => q_4_0_54_port, B => q_4_1_54_port, Ci =>
                           q_4_2_54_port, S => q_5_0_54_port, Co => 
                           q_5_1_55_port);
   FA_C_4_0_55 : FA_195 port map( A => q_4_0_55_port, B => q_4_1_55_port, Ci =>
                           q_4_2_55_port, S => q_5_0_55_port, Co => 
                           q_5_1_56_port);
   FA_C_4_0_56 : FA_194 port map( A => q_4_0_56_port, B => q_4_1_56_port, Ci =>
                           q_4_2_56_port, S => q_5_0_56_port, Co => 
                           q_5_1_57_port);
   FA_C_4_0_57 : FA_193 port map( A => q_4_0_57_port, B => q_4_1_57_port, Ci =>
                           q_4_2_57_port, S => q_5_0_57_port, Co => 
                           q_5_1_58_port);
   FA_C_4_0_58 : FA_192 port map( A => q_4_0_58_port, B => q_4_1_58_port, Ci =>
                           q_4_2_58_port, S => q_5_0_58_port, Co => 
                           q_5_1_59_port);
   FA_C_4_0_59 : FA_191 port map( A => q_4_0_59_port, B => q_4_1_59_port, Ci =>
                           q_4_2_59_port, S => q_5_0_59_port, Co => 
                           q_5_1_60_port);
   FA_C_4_0_60 : FA_190 port map( A => q_4_0_60_port, B => q_4_1_60_port, Ci =>
                           q_0_2_60_port, S => q_5_0_60_port, Co => 
                           q_5_1_61_port);
   FA_C_4_0_61 : FA_189 port map( A => q_4_0_61_port, B => n82, Ci => 
                           q_0_1_61_port, S => q_5_0_61_port, Co => 
                           q_5_1_62_port);
   HA_L_4_0_62 : HA_3 port map( A => X_Logic1_port, B => q_0_1_62_port, S => 
                           q_5_0_62_port, C => q_5_0_63_port);
   HA_R_5_0_2 : HA_2 port map( A => q_0_0_2_port, B => q_0_1_2_port, S => 
                           q_6_0_2_port, C => q_6_1_3_port);
   HA_R_5_0_3 : HA_1 port map( A => q_0_0_3_port, B => q_0_1_3_port, S => 
                           q_6_0_3_port, C => q_6_1_4_port);
   FA_C_5_0_4 : FA_188 port map( A => q_5_0_4_port, B => q_0_2_4_port, Ci => 
                           n10, S => q_6_0_4_port, Co => q_6_1_5_port);
   FA_C_5_0_5 : FA_187 port map( A => q_5_0_5_port, B => q_5_1_5_port, Ci => 
                           q_0_2_5_port, S => q_6_0_5_port, Co => q_6_1_6_port)
                           ;
   FA_C_5_0_6 : FA_186 port map( A => q_5_0_6_port, B => q_5_1_6_port, Ci => 
                           n14, S => q_6_0_6_port, Co => q_6_1_7_port);
   FA_C_5_0_7 : FA_185 port map( A => q_5_0_7_port, B => q_5_1_7_port, Ci => 
                           q_0_3_7_port, S => q_6_0_7_port, Co => q_6_1_8_port)
                           ;
   FA_C_5_0_8 : FA_184 port map( A => q_5_0_8_port, B => q_5_1_8_port, Ci => n8
                           , S => q_6_0_8_port, Co => q_6_1_9_port);
   FA_C_5_0_9 : FA_183 port map( A => q_5_0_9_port, B => q_5_1_9_port, Ci => 
                           q_5_2_9_port, S => q_6_0_9_port, Co => q_6_1_10_port
                           );
   FA_C_5_0_10 : FA_182 port map( A => q_5_0_10_port, B => q_5_1_10_port, Ci =>
                           q_5_2_10_port, S => q_6_0_10_port, Co => 
                           q_6_1_11_port);
   FA_C_5_0_11 : FA_181 port map( A => q_5_0_11_port, B => q_5_1_11_port, Ci =>
                           q_5_2_11_port, S => q_6_0_11_port, Co => 
                           q_6_1_12_port);
   FA_C_5_0_12 : FA_180 port map( A => q_5_0_12_port, B => q_5_1_12_port, Ci =>
                           q_5_2_12_port, S => q_6_0_12_port, Co => 
                           q_6_1_13_port);
   FA_C_5_0_13 : FA_179 port map( A => q_5_0_13_port, B => q_5_1_13_port, Ci =>
                           q_5_2_13_port, S => q_6_0_13_port, Co => 
                           q_6_1_14_port);
   FA_C_5_0_14 : FA_178 port map( A => q_5_0_14_port, B => q_5_1_14_port, Ci =>
                           q_5_2_14_port, S => q_6_0_14_port, Co => 
                           q_6_1_15_port);
   FA_C_5_0_15 : FA_177 port map( A => q_5_0_15_port, B => q_5_1_15_port, Ci =>
                           q_5_2_15_port, S => q_6_0_15_port, Co => 
                           q_6_1_16_port);
   FA_C_5_0_16 : FA_176 port map( A => q_5_0_16_port, B => q_5_1_16_port, Ci =>
                           q_5_2_16_port, S => q_6_0_16_port, Co => 
                           q_6_1_17_port);
   FA_C_5_0_17 : FA_175 port map( A => q_5_0_17_port, B => q_5_1_17_port, Ci =>
                           q_5_2_17_port, S => q_6_0_17_port, Co => 
                           q_6_1_18_port);
   FA_C_5_0_18 : FA_174 port map( A => q_5_0_18_port, B => q_5_1_18_port, Ci =>
                           q_5_2_18_port, S => q_6_0_18_port, Co => 
                           q_6_1_19_port);
   FA_C_5_0_19 : FA_173 port map( A => q_5_0_19_port, B => q_5_1_19_port, Ci =>
                           q_5_2_19_port, S => q_6_0_19_port, Co => 
                           q_6_1_20_port);
   FA_C_5_0_20 : FA_172 port map( A => q_5_0_20_port, B => q_5_1_20_port, Ci =>
                           q_5_2_20_port, S => q_6_0_20_port, Co => 
                           q_6_1_21_port);
   FA_C_5_0_21 : FA_171 port map( A => q_5_0_21_port, B => q_5_1_21_port, Ci =>
                           q_5_2_21_port, S => q_6_0_21_port, Co => 
                           q_6_1_22_port);
   FA_C_5_0_22 : FA_170 port map( A => q_5_0_22_port, B => q_5_1_22_port, Ci =>
                           q_5_2_22_port, S => q_6_0_22_port, Co => 
                           q_6_1_23_port);
   FA_C_5_0_23 : FA_169 port map( A => q_5_0_23_port, B => q_5_1_23_port, Ci =>
                           q_5_2_23_port, S => q_6_0_23_port, Co => 
                           q_6_1_24_port);
   FA_C_5_0_24 : FA_168 port map( A => q_5_0_24_port, B => q_5_1_24_port, Ci =>
                           q_5_2_24_port, S => q_6_0_24_port, Co => 
                           q_6_1_25_port);
   FA_C_5_0_25 : FA_167 port map( A => q_5_0_25_port, B => q_5_1_25_port, Ci =>
                           q_5_2_25_port, S => q_6_0_25_port, Co => 
                           q_6_1_26_port);
   FA_C_5_0_26 : FA_166 port map( A => q_5_0_26_port, B => q_5_1_26_port, Ci =>
                           q_5_2_26_port, S => q_6_0_26_port, Co => 
                           q_6_1_27_port);
   FA_C_5_0_27 : FA_165 port map( A => q_5_0_27_port, B => q_5_1_27_port, Ci =>
                           q_5_2_27_port, S => q_6_0_27_port, Co => 
                           q_6_1_28_port);
   FA_C_5_0_28 : FA_164 port map( A => q_5_0_28_port, B => q_5_1_28_port, Ci =>
                           q_5_2_28_port, S => q_6_0_28_port, Co => 
                           q_6_1_29_port);
   FA_C_5_0_29 : FA_163 port map( A => q_5_0_29_port, B => q_5_1_29_port, Ci =>
                           q_5_2_29_port, S => q_6_0_29_port, Co => 
                           q_6_1_30_port);
   FA_C_5_0_30 : FA_162 port map( A => q_5_0_30_port, B => q_5_1_30_port, Ci =>
                           q_5_2_30_port, S => q_6_0_30_port, Co => 
                           q_6_1_31_port);
   FA_C_5_0_31 : FA_161 port map( A => q_5_0_31_port, B => q_5_1_31_port, Ci =>
                           q_5_2_31_port, S => q_6_0_31_port, Co => 
                           q_6_1_32_port);
   FA_C_5_0_32 : FA_160 port map( A => q_5_0_32_port, B => q_5_1_32_port, Ci =>
                           q_5_2_32_port, S => q_6_0_32_port, Co => 
                           q_6_1_33_port);
   FA_C_5_0_33 : FA_159 port map( A => q_5_0_33_port, B => q_5_1_33_port, Ci =>
                           q_5_2_33_port, S => q_6_0_33_port, Co => 
                           q_6_1_34_port);
   FA_C_5_0_34 : FA_158 port map( A => q_5_0_34_port, B => q_5_1_34_port, Ci =>
                           q_5_2_34_port, S => q_6_0_34_port, Co => 
                           q_6_1_35_port);
   FA_C_5_0_35 : FA_157 port map( A => q_5_0_35_port, B => q_5_1_35_port, Ci =>
                           q_5_2_35_port, S => q_6_0_35_port, Co => 
                           q_6_1_36_port);
   FA_C_5_0_36 : FA_156 port map( A => q_5_0_36_port, B => q_5_1_36_port, Ci =>
                           q_5_2_36_port, S => q_6_0_36_port, Co => 
                           q_6_1_37_port);
   FA_C_5_0_37 : FA_155 port map( A => q_5_0_37_port, B => q_5_1_37_port, Ci =>
                           q_5_2_37_port, S => q_6_0_37_port, Co => 
                           q_6_1_38_port);
   FA_C_5_0_38 : FA_154 port map( A => q_5_0_38_port, B => q_5_1_38_port, Ci =>
                           q_5_2_38_port, S => q_6_0_38_port, Co => 
                           q_6_1_39_port);
   FA_C_5_0_39 : FA_153 port map( A => q_5_0_39_port, B => q_5_1_39_port, Ci =>
                           q_5_2_39_port, S => q_6_0_39_port, Co => 
                           q_6_1_40_port);
   FA_C_5_0_40 : FA_152 port map( A => q_5_0_40_port, B => q_5_1_40_port, Ci =>
                           q_5_2_40_port, S => q_6_0_40_port, Co => 
                           q_6_1_41_port);
   FA_C_5_0_41 : FA_151 port map( A => q_5_0_41_port, B => q_5_1_41_port, Ci =>
                           q_5_2_41_port, S => q_6_0_41_port, Co => 
                           q_6_1_42_port);
   FA_C_5_0_42 : FA_150 port map( A => q_5_0_42_port, B => q_5_1_42_port, Ci =>
                           q_5_2_42_port, S => q_6_0_42_port, Co => 
                           q_6_1_43_port);
   FA_C_5_0_43 : FA_149 port map( A => q_5_0_43_port, B => q_5_1_43_port, Ci =>
                           q_5_2_43_port, S => q_6_0_43_port, Co => 
                           q_6_1_44_port);
   FA_C_5_0_44 : FA_148 port map( A => q_5_0_44_port, B => q_5_1_44_port, Ci =>
                           q_5_2_44_port, S => q_6_0_44_port, Co => 
                           q_6_1_45_port);
   FA_C_5_0_45 : FA_147 port map( A => q_5_0_45_port, B => q_5_1_45_port, Ci =>
                           q_5_2_45_port, S => q_6_0_45_port, Co => 
                           q_6_1_46_port);
   FA_C_5_0_46 : FA_146 port map( A => q_5_0_46_port, B => q_5_1_46_port, Ci =>
                           q_5_2_46_port, S => q_6_0_46_port, Co => 
                           q_6_1_47_port);
   FA_C_5_0_47 : FA_145 port map( A => q_5_0_47_port, B => q_5_1_47_port, Ci =>
                           q_5_2_47_port, S => q_6_0_47_port, Co => 
                           q_6_1_48_port);
   FA_C_5_0_48 : FA_144 port map( A => q_5_0_48_port, B => q_5_1_48_port, Ci =>
                           q_5_2_48_port, S => q_6_0_48_port, Co => 
                           q_6_1_49_port);
   FA_C_5_0_49 : FA_143 port map( A => q_5_0_49_port, B => q_5_1_49_port, Ci =>
                           q_5_2_49_port, S => q_6_0_49_port, Co => 
                           q_6_1_50_port);
   FA_C_5_0_50 : FA_142 port map( A => q_5_0_50_port, B => q_5_1_50_port, Ci =>
                           q_5_2_50_port, S => q_6_0_50_port, Co => 
                           q_6_1_51_port);
   FA_C_5_0_51 : FA_141 port map( A => q_5_0_51_port, B => q_5_1_51_port, Ci =>
                           q_5_2_51_port, S => q_6_0_51_port, Co => 
                           q_6_1_52_port);
   FA_C_5_0_52 : FA_140 port map( A => q_5_0_52_port, B => q_5_1_52_port, Ci =>
                           q_5_2_52_port, S => q_6_0_52_port, Co => 
                           q_6_1_53_port);
   FA_C_5_0_53 : FA_139 port map( A => q_5_0_53_port, B => q_5_1_53_port, Ci =>
                           q_5_2_53_port, S => q_6_0_53_port, Co => 
                           q_6_1_54_port);
   FA_C_5_0_54 : FA_138 port map( A => q_5_0_54_port, B => q_5_1_54_port, Ci =>
                           q_5_2_54_port, S => q_6_0_54_port, Co => 
                           q_6_1_55_port);
   FA_C_5_0_55 : FA_137 port map( A => q_5_0_55_port, B => q_5_1_55_port, Ci =>
                           q_5_2_55_port, S => q_6_0_55_port, Co => 
                           q_6_1_56_port);
   FA_C_5_0_56 : FA_136 port map( A => q_5_0_56_port, B => q_5_1_56_port, Ci =>
                           q_5_2_56_port, S => q_6_0_56_port, Co => 
                           q_6_1_57_port);
   FA_C_5_0_57 : FA_135 port map( A => q_5_0_57_port, B => q_5_1_57_port, Ci =>
                           q_5_2_57_port, S => q_6_0_57_port, Co => 
                           q_6_1_58_port);
   FA_C_5_0_58 : FA_134 port map( A => q_5_0_58_port, B => q_5_1_58_port, Ci =>
                           q_5_2_58_port, S => q_6_0_58_port, Co => 
                           q_6_1_59_port);
   FA_C_5_0_59 : FA_133 port map( A => q_5_0_59_port, B => q_5_1_59_port, Ci =>
                           q_0_3_59_port, S => q_6_0_59_port, Co => 
                           q_6_1_60_port);
   FA_C_5_0_60 : FA_132 port map( A => q_5_0_60_port, B => q_5_1_60_port, Ci =>
                           q_0_3_60_port, S => q_6_0_60_port, Co => 
                           q_6_1_61_port);
   FA_C_5_0_61 : FA_131 port map( A => q_5_0_61_port, B => q_5_1_61_port, Ci =>
                           q_0_2_61_port, S => q_6_0_61_port, Co => 
                           q_6_1_62_port);
   FA_C_5_0_62 : FA_130 port map( A => q_5_0_62_port, B => q_5_1_62_port, Ci =>
                           q_0_2_62_port, S => q_6_0_62_port, Co => 
                           q_6_1_63_port);
   FA_C_5_5_0_63 : FA_129 port map( A => q_5_0_63_port, B => n81, Ci => 
                           q_0_1_63_port, S => q_6_0_63_port, Co => n_1043);
   P4_ADDER_0 : P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16 port map( A(63) => 
                           q_6_0_63_port, A(62) => q_6_0_62_port, A(61) => 
                           q_6_0_61_port, A(60) => q_6_0_60_port, A(59) => 
                           q_6_0_59_port, A(58) => q_6_0_58_port, A(57) => 
                           q_6_0_57_port, A(56) => q_6_0_56_port, A(55) => 
                           q_6_0_55_port, A(54) => q_6_0_54_port, A(53) => 
                           q_6_0_53_port, A(52) => q_6_0_52_port, A(51) => 
                           q_6_0_51_port, A(50) => q_6_0_50_port, A(49) => 
                           q_6_0_49_port, A(48) => q_6_0_48_port, A(47) => 
                           q_6_0_47_port, A(46) => q_6_0_46_port, A(45) => 
                           q_6_0_45_port, A(44) => q_6_0_44_port, A(43) => 
                           q_6_0_43_port, A(42) => q_6_0_42_port, A(41) => 
                           q_6_0_41_port, A(40) => q_6_0_40_port, A(39) => 
                           q_6_0_39_port, A(38) => q_6_0_38_port, A(37) => 
                           q_6_0_37_port, A(36) => q_6_0_36_port, A(35) => 
                           q_6_0_35_port, A(34) => q_6_0_34_port, A(33) => 
                           q_6_0_33_port, A(32) => q_6_0_32_port, A(31) => 
                           q_6_0_31_port, A(30) => q_6_0_30_port, A(29) => 
                           q_6_0_29_port, A(28) => q_6_0_28_port, A(27) => 
                           q_6_0_27_port, A(26) => q_6_0_26_port, A(25) => 
                           q_6_0_25_port, A(24) => q_6_0_24_port, A(23) => 
                           q_6_0_23_port, A(22) => q_6_0_22_port, A(21) => 
                           q_6_0_21_port, A(20) => q_6_0_20_port, A(19) => 
                           q_6_0_19_port, A(18) => q_6_0_18_port, A(17) => 
                           q_6_0_17_port, A(16) => q_6_0_16_port, A(15) => 
                           q_6_0_15_port, A(14) => q_6_0_14_port, A(13) => 
                           q_6_0_13_port, A(12) => q_6_0_12_port, A(11) => 
                           q_6_0_11_port, A(10) => q_6_0_10_port, A(9) => 
                           q_6_0_9_port, A(8) => q_6_0_8_port, A(7) => 
                           q_6_0_7_port, A(6) => q_6_0_6_port, A(5) => 
                           q_6_0_5_port, A(4) => q_6_0_4_port, A(3) => 
                           q_6_0_3_port, A(2) => q_6_0_2_port, A(1) => 
                           q_0_0_1_port, A(0) => q_0_0_0_port, B(63) => 
                           q_6_1_63_port, B(62) => q_6_1_62_port, B(61) => 
                           q_6_1_61_port, B(60) => q_6_1_60_port, B(59) => 
                           q_6_1_59_port, B(58) => q_6_1_58_port, B(57) => 
                           q_6_1_57_port, B(56) => q_6_1_56_port, B(55) => 
                           q_6_1_55_port, B(54) => q_6_1_54_port, B(53) => 
                           q_6_1_53_port, B(52) => q_6_1_52_port, B(51) => 
                           q_6_1_51_port, B(50) => q_6_1_50_port, B(49) => 
                           q_6_1_49_port, B(48) => q_6_1_48_port, B(47) => 
                           q_6_1_47_port, B(46) => q_6_1_46_port, B(45) => 
                           q_6_1_45_port, B(44) => q_6_1_44_port, B(43) => 
                           q_6_1_43_port, B(42) => q_6_1_42_port, B(41) => 
                           q_6_1_41_port, B(40) => q_6_1_40_port, B(39) => 
                           q_6_1_39_port, B(38) => q_6_1_38_port, B(37) => 
                           q_6_1_37_port, B(36) => q_6_1_36_port, B(35) => 
                           q_6_1_35_port, B(34) => q_6_1_34_port, B(33) => 
                           q_6_1_33_port, B(32) => q_6_1_32_port, B(31) => 
                           q_6_1_31_port, B(30) => q_6_1_30_port, B(29) => 
                           q_6_1_29_port, B(28) => q_6_1_28_port, B(27) => 
                           q_6_1_27_port, B(26) => q_6_1_26_port, B(25) => 
                           q_6_1_25_port, B(24) => q_6_1_24_port, B(23) => 
                           q_6_1_23_port, B(22) => q_6_1_22_port, B(21) => 
                           q_6_1_21_port, B(20) => q_6_1_20_port, B(19) => 
                           q_6_1_19_port, B(18) => q_6_1_18_port, B(17) => 
                           q_6_1_17_port, B(16) => q_6_1_16_port, B(15) => 
                           q_6_1_15_port, B(14) => q_6_1_14_port, B(13) => 
                           q_6_1_13_port, B(12) => q_6_1_12_port, B(11) => 
                           q_6_1_11_port, B(10) => q_6_1_10_port, B(9) => 
                           q_6_1_9_port, B(8) => q_6_1_8_port, B(7) => 
                           q_6_1_7_port, B(6) => q_6_1_6_port, B(5) => 
                           q_6_1_5_port, B(4) => q_6_1_4_port, B(3) => 
                           q_6_1_3_port, B(2) => n16, B(1) => X_Logic0_port, 
                           B(0) => n15, Cin => X_Logic0_port, S(63) => C(63), 
                           S(62) => C(62), S(61) => C(61), S(60) => C(60), 
                           S(59) => C(59), S(58) => C(58), S(57) => C(57), 
                           S(56) => C(56), S(55) => C(55), S(54) => C(54), 
                           S(53) => C(53), S(52) => C(52), S(51) => C(51), 
                           S(50) => C(50), S(49) => C(49), S(48) => C(48), 
                           S(47) => C(47), S(46) => C(46), S(45) => C(45), 
                           S(44) => C(44), S(43) => C(43), S(42) => C(42), 
                           S(41) => C(41), S(40) => C(40), S(39) => C(39), 
                           S(38) => C(38), S(37) => C(37), S(36) => C(36), 
                           S(35) => C(35), S(34) => C(34), S(33) => C(33), 
                           S(32) => C(32), S(31) => C(31), S(30) => C(30), 
                           S(29) => C(29), S(28) => C(28), S(27) => C(27), 
                           S(26) => C(26), S(25) => C(25), S(24) => C(24), 
                           S(23) => C(23), S(22) => C(22), S(21) => C(21), 
                           S(20) => C(20), S(19) => C(19), S(18) => C(18), 
                           S(17) => C(17), S(16) => C(16), S(15) => C(15), 
                           S(14) => C(14), S(13) => C(13), S(12) => C(12), 
                           S(11) => C(11), S(10) => C(10), S(9) => C(9), S(8) 
                           => C(8), S(7) => C(7), S(6) => C(6), S(5) => C(5), 
                           S(4) => C(4), S(3) => C(3), S(2) => C(2), S(1) => 
                           C(1), S(0) => C(0), Cout => n_1044);
   U3 : CLKBUF_X1 port map( A => B(13), Z => n1);
   U4 : CLKBUF_X1 port map( A => B(1), Z => n2);
   U5 : BUF_X2 port map( A => B(23), Z => n3);
   U6 : CLKBUF_X1 port map( A => B(21), Z => n4);
   U7 : CLKBUF_X1 port map( A => B(11), Z => n5);
   U8 : BUF_X4 port map( A => A(21), Z => n60);
   U9 : CLKBUF_X1 port map( A => n3, Z => n6);
   U10 : CLKBUF_X1 port map( A => B(17), Z => n7);
   U11 : CLKBUF_X1 port map( A => B(9), Z => n8);
   U12 : CLKBUF_X1 port map( A => B(19), Z => n9);
   U13 : CLKBUF_X1 port map( A => B(5), Z => n10);
   U14 : CLKBUF_X1 port map( A => B(7), Z => n11);
   U15 : CLKBUF_X1 port map( A => n2, Z => n12);
   U16 : CLKBUF_X1 port map( A => B(15), Z => n13);
   U17 : CLKBUF_X1 port map( A => n11, Z => n14);
   U18 : CLKBUF_X3 port map( A => A(10), Z => n37);
   U19 : CLKBUF_X1 port map( A => A(1), Z => n20);
   U20 : CLKBUF_X1 port map( A => A(4), Z => n26);
   U21 : CLKBUF_X3 port map( A => A(7), Z => n31);
   U22 : CLKBUF_X1 port map( A => A(6), Z => n30);
   U23 : CLKBUF_X1 port map( A => A(5), Z => n28);
   U24 : BUF_X4 port map( A => A(1), Z => n19);
   U25 : BUF_X4 port map( A => A(4), Z => n25);
   U26 : BUF_X4 port map( A => A(9), Z => n35);
   U27 : CLKBUF_X1 port map( A => B(3), Z => n16);
   U28 : INV_X1 port map( A => n96, ZN => n15);
   U29 : CLKBUF_X3 port map( A => A(14), Z => n45);
   U30 : CLKBUF_X3 port map( A => A(2), Z => n21);
   U31 : CLKBUF_X3 port map( A => A(3), Z => n23);
   U32 : CLKBUF_X3 port map( A => A(15), Z => n47);
   U33 : CLKBUF_X3 port map( A => A(17), Z => n51);
   U34 : CLKBUF_X3 port map( A => A(0), Z => n17);
   U35 : CLKBUF_X3 port map( A => A(5), Z => n27);
   U36 : CLKBUF_X3 port map( A => A(6), Z => n29);
   U37 : CLKBUF_X3 port map( A => A(8), Z => n33);
   U38 : CLKBUF_X3 port map( A => A(23), Z => n63);
   U39 : CLKBUF_X3 port map( A => A(11), Z => n39);
   U40 : CLKBUF_X3 port map( A => A(12), Z => n41);
   U41 : CLKBUF_X3 port map( A => A(13), Z => n43);
   U42 : CLKBUF_X3 port map( A => A(22), Z => n61);
   U43 : CLKBUF_X3 port map( A => A(19), Z => n55);
   U44 : CLKBUF_X3 port map( A => A(16), Z => n49);
   U45 : CLKBUF_X3 port map( A => A(20), Z => n57);
   U46 : CLKBUF_X3 port map( A => A(18), Z => n53);
   U47 : BUF_X1 port map( A => A(10), Z => n38);
   U48 : BUF_X1 port map( A => A(9), Z => n36);
   U49 : BUF_X1 port map( A => A(14), Z => n46);
   U50 : BUF_X1 port map( A => A(13), Z => n44);
   U51 : BUF_X1 port map( A => A(11), Z => n40);
   U52 : BUF_X1 port map( A => A(7), Z => n32);
   U53 : BUF_X1 port map( A => A(12), Z => n42);
   U54 : BUF_X1 port map( A => A(8), Z => n34);
   U55 : CLKBUF_X1 port map( A => A(3), Z => n24);
   U56 : CLKBUF_X1 port map( A => A(2), Z => n22);
   U57 : CLKBUF_X1 port map( A => A(0), Z => n18);
   U58 : BUF_X2 port map( A => A(16), Z => n50);
   U59 : BUF_X2 port map( A => A(15), Z => n48);
   U60 : BUF_X2 port map( A => A(18), Z => n54);
   U61 : BUF_X2 port map( A => A(17), Z => n52);
   U62 : BUF_X1 port map( A => A(20), Z => n58);
   U63 : BUF_X1 port map( A => A(19), Z => n56);
   U64 : BUF_X2 port map( A => A(22), Z => n62);
   U65 : CLKBUF_X1 port map( A => A(23), Z => n64);
   U66 : INV_X1 port map( A => n6, ZN => n85);
   U67 : INV_X1 port map( A => n4, ZN => n86);
   U68 : INV_X1 port map( A => n9, ZN => n87);
   U69 : INV_X1 port map( A => n7, ZN => n88);
   U70 : BUF_X2 port map( A => A(24), Z => n65);
   U71 : BUF_X2 port map( A => A(25), Z => n67);
   U72 : BUF_X2 port map( A => A(26), Z => n69);
   U73 : BUF_X2 port map( A => A(28), Z => n73);
   U74 : BUF_X2 port map( A => A(27), Z => n71);
   U75 : BUF_X2 port map( A => A(29), Z => n75);
   U76 : BUF_X2 port map( A => A(30), Z => n77);
   U77 : BUF_X1 port map( A => A(25), Z => n68);
   U78 : BUF_X1 port map( A => A(29), Z => n76);
   U79 : BUF_X1 port map( A => A(24), Z => n66);
   U80 : BUF_X1 port map( A => A(26), Z => n70);
   U81 : BUF_X1 port map( A => A(30), Z => n78);
   U82 : BUF_X1 port map( A => A(27), Z => n72);
   U83 : BUF_X1 port map( A => A(28), Z => n74);
   U84 : BUF_X1 port map( A => A(31), Z => n80);
   U85 : INV_X1 port map( A => B(27), ZN => n83);
   U86 : INV_X1 port map( A => B(25), ZN => n84);
   U87 : INV_X1 port map( A => B(29), ZN => n82);
   U88 : INV_X1 port map( A => B(31), ZN => n81);
   U89 : CLKBUF_X1 port map( A => A(21), Z => n59);
   U90 : CLKBUF_X1 port map( A => A(31), Z => n79);
   U91 : INV_X1 port map( A => B(15), ZN => n89);
   U92 : INV_X1 port map( A => n1, ZN => n90);
   U93 : INV_X1 port map( A => n5, ZN => n91);
   U94 : INV_X1 port map( A => n8, ZN => n92);
   U95 : INV_X1 port map( A => n11, ZN => n93);
   U96 : INV_X1 port map( A => n10, ZN => n94);
   U97 : INV_X1 port map( A => n16, ZN => n95);
   U98 : INV_X1 port map( A => n2, ZN => n96);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity UnpackFP_0 is

   port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector 
         (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, isNaN,
         isINF, isZ, isDN : out std_logic);

end UnpackFP_0;

architecture SYN_UnpackFP of UnpackFP_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, N13, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12
      , n13_port, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, 
      n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37 : std_logic;

begin
   SIG <= ( X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, 
      X_Logic0_port, X_Logic0_port, X_Logic0_port, X_Logic0_port, N13, FP(22), 
      FP(21), FP(20), FP(19), FP(18), FP(17), FP(16), FP(15), FP(14), FP(13), 
      FP(12), FP(11), FP(10), FP(9), FP(8), FP(7), FP(6), FP(5), FP(4), FP(3), 
      FP(2), FP(1), FP(0) );
   EXP <= ( FP(30), FP(29), FP(28), FP(27), FP(26), FP(25), FP(24), FP(23) );
   SIGN <= FP(31);
   
   X_Logic0_port <= '0';
   U2 : NAND4_X1 port map( A1 => n24, A2 => n23, A3 => n22, A4 => n21, ZN => 
                           n35);
   U3 : NOR2_X1 port map( A1 => FP(0), A2 => FP(1), ZN => n24);
   U4 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => n22);
   U5 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U6 : NOR2_X1 port map( A1 => FP(10), A2 => FP(9), ZN => n3);
   U7 : INV_X1 port map( A => FP(19), ZN => n17);
   U8 : INV_X1 port map( A => FP(20), ZN => n16);
   U9 : NOR2_X1 port map( A1 => FP(18), A2 => FP(17), ZN => n18);
   U10 : INV_X1 port map( A => FP(13), ZN => n12);
   U11 : INV_X1 port map( A => FP(14), ZN => n11);
   U12 : NOR2_X1 port map( A1 => FP(12), A2 => FP(11), ZN => n13_port);
   U13 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n23);
   U14 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n9);
   U15 : NAND4_X1 port map( A1 => n6, A2 => n5, A3 => n4, A4 => n3, ZN => n10);
   U16 : INV_X1 port map( A => FP(4), ZN => n7);
   U17 : NOR2_X1 port map( A1 => FP(3), A2 => FP(2), ZN => n8);
   U18 : NOR2_X1 port map( A1 => FP(5), A2 => FP(6), ZN => n6);
   U19 : OR2_X1 port map( A1 => FP(22), A2 => FP(21), ZN => n19);
   U20 : OR2_X1 port map( A1 => FP(16), A2 => FP(15), ZN => n14);
   U21 : INV_X1 port map( A => FP(8), ZN => n4);
   U22 : INV_X1 port map( A => FP(7), ZN => n5);
   U23 : NOR4_X1 port map( A1 => FP(27), A2 => FP(28), A3 => FP(29), A4 => 
                           FP(30), ZN => n2);
   U24 : NOR4_X1 port map( A1 => FP(23), A2 => FP(24), A3 => FP(25), A4 => 
                           FP(26), ZN => n1);
   U25 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => N13);
   U26 : NAND3_X1 port map( A1 => n13_port, A2 => n12, A3 => n11, ZN => n15);
   U27 : NAND3_X1 port map( A1 => n18, A2 => n17, A3 => n16, ZN => n20);
   U28 : INV_X1 port map( A => n35, ZN => n37);
   U29 : NOR2_X1 port map( A1 => N13, A2 => n37, ZN => isDN);
   U30 : NOR2_X1 port map( A1 => N13, A2 => n35, ZN => isZ);
   U31 : INV_X1 port map( A => FP(28), ZN => n28);
   U32 : INV_X1 port map( A => FP(27), ZN => n27);
   U33 : INV_X1 port map( A => FP(30), ZN => n26);
   U34 : INV_X1 port map( A => FP(29), ZN => n25);
   U35 : NOR4_X1 port map( A1 => n28, A2 => n27, A3 => n26, A4 => n25, ZN => 
                           n34);
   U36 : INV_X1 port map( A => FP(24), ZN => n32);
   U37 : INV_X1 port map( A => FP(23), ZN => n31);
   U38 : INV_X1 port map( A => FP(26), ZN => n30);
   U39 : INV_X1 port map( A => FP(25), ZN => n29);
   U40 : NOR4_X1 port map( A1 => n32, A2 => n31, A3 => n30, A4 => n29, ZN => 
                           n33);
   U41 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => n36);
   U42 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => isINF);
   U43 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => isNaN);

end SYN_UnpackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage4 is

   port( EXP_neg : in std_logic;  EXP_out_round : in std_logic_vector (7 downto
         0);  EXP_pos, SIGN_out : in std_logic;  SIG_out_round : in 
         std_logic_vector (27 downto 0);  clk, isINF_tab, isNaN, isZ_tab : in 
         std_logic;  FP_Z : out std_logic_vector (31 downto 0));

end FPmul_stage4;

architecture SYN_struct of FPmul_stage4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component PackFP
      port( SIGN : in std_logic;  EXP : in std_logic_vector (7 downto 0);  SIG 
            : in std_logic_vector (22 downto 0);  isNaN, isINF, isZ : in 
            std_logic;  FP : out std_logic_vector (31 downto 0));
   end component;
   
   component FPnormalize_SIG_width28_1
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0));
   end component;
   
   signal SIG_out_norm2_26_port, SIG_out_22_port, SIG_out_21_port, 
      SIG_out_20_port, SIG_out_19_port, SIG_out_18_port, SIG_out_17_port, 
      SIG_out_16_port, SIG_out_15_port, SIG_out_14_port, SIG_out_13_port, 
      SIG_out_12_port, SIG_out_11_port, SIG_out_10_port, SIG_out_9_port, 
      SIG_out_8_port, SIG_out_7_port, SIG_out_6_port, SIG_out_5_port, 
      SIG_out_4_port, SIG_out_3_port, SIG_out_2_port, SIG_out_1_port, 
      SIG_out_0_port, EXP_out_7_port, EXP_out_6_port, EXP_out_5_port, 
      EXP_out_4_port, EXP_out_3_port, EXP_out_2_port, EXP_out_1_port, 
      EXP_out_0_port, isINF, FP_31_port, FP_30_port, FP_29_port, FP_28_port, 
      FP_27_port, FP_26_port, FP_25_port, FP_24_port, FP_23_port, FP_22_port, 
      FP_21_port, FP_20_port, FP_19_port, FP_18_port, FP_17_port, FP_16_port, 
      FP_15_port, FP_14_port, FP_13_port, FP_12_port, FP_11_port, FP_10_port, 
      FP_9_port, FP_8_port, FP_7_port, FP_6_port, FP_5_port, FP_4_port, 
      FP_3_port, FP_2_port, FP_1_port, FP_0_port, n1, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, 
      n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, 
      n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, 
      n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080 : std_logic;

begin
   
   I1 : FPnormalize_SIG_width28_1 port map( SIG_in(27) => SIG_out_round(27), 
                           SIG_in(26) => SIG_out_round(26), SIG_in(25) => 
                           SIG_out_round(25), SIG_in(24) => SIG_out_round(24), 
                           SIG_in(23) => SIG_out_round(23), SIG_in(22) => 
                           SIG_out_round(22), SIG_in(21) => SIG_out_round(21), 
                           SIG_in(20) => SIG_out_round(20), SIG_in(19) => 
                           SIG_out_round(19), SIG_in(18) => SIG_out_round(18), 
                           SIG_in(17) => SIG_out_round(17), SIG_in(16) => 
                           SIG_out_round(16), SIG_in(15) => SIG_out_round(15), 
                           SIG_in(14) => SIG_out_round(14), SIG_in(13) => 
                           SIG_out_round(13), SIG_in(12) => SIG_out_round(12), 
                           SIG_in(11) => SIG_out_round(11), SIG_in(10) => 
                           SIG_out_round(10), SIG_in(9) => SIG_out_round(9), 
                           SIG_in(8) => SIG_out_round(8), SIG_in(7) => 
                           SIG_out_round(7), SIG_in(6) => SIG_out_round(6), 
                           SIG_in(5) => SIG_out_round(5), SIG_in(4) => 
                           SIG_out_round(4), SIG_in(3) => SIG_out_round(3), 
                           SIG_in(2) => SIG_out_round(2), SIG_in(1) => 
                           SIG_out_round(1), SIG_in(0) => SIG_out_round(0), 
                           EXP_in(7) => EXP_out_round(7), EXP_in(6) => 
                           EXP_out_round(6), EXP_in(5) => EXP_out_round(5), 
                           EXP_in(4) => EXP_out_round(4), EXP_in(3) => 
                           EXP_out_round(3), EXP_in(2) => EXP_out_round(2), 
                           EXP_in(1) => EXP_out_round(1), EXP_in(0) => 
                           EXP_out_round(0), SIG_out(27) => n_1045, SIG_out(26)
                           => SIG_out_norm2_26_port, SIG_out(25) => 
                           SIG_out_22_port, SIG_out(24) => SIG_out_21_port, 
                           SIG_out(23) => SIG_out_20_port, SIG_out(22) => 
                           SIG_out_19_port, SIG_out(21) => SIG_out_18_port, 
                           SIG_out(20) => SIG_out_17_port, SIG_out(19) => 
                           SIG_out_16_port, SIG_out(18) => SIG_out_15_port, 
                           SIG_out(17) => SIG_out_14_port, SIG_out(16) => 
                           SIG_out_13_port, SIG_out(15) => SIG_out_12_port, 
                           SIG_out(14) => SIG_out_11_port, SIG_out(13) => 
                           SIG_out_10_port, SIG_out(12) => SIG_out_9_port, 
                           SIG_out(11) => SIG_out_8_port, SIG_out(10) => 
                           SIG_out_7_port, SIG_out(9) => SIG_out_6_port, 
                           SIG_out(8) => SIG_out_5_port, SIG_out(7) => 
                           SIG_out_4_port, SIG_out(6) => SIG_out_3_port, 
                           SIG_out(5) => SIG_out_2_port, SIG_out(4) => 
                           SIG_out_1_port, SIG_out(3) => SIG_out_0_port, 
                           SIG_out(2) => n_1046, SIG_out(1) => n_1047, 
                           SIG_out(0) => n_1048, EXP_out(7) => EXP_out_7_port, 
                           EXP_out(6) => EXP_out_6_port, EXP_out(5) => 
                           EXP_out_5_port, EXP_out(4) => EXP_out_4_port, 
                           EXP_out(3) => EXP_out_3_port, EXP_out(2) => 
                           EXP_out_2_port, EXP_out(1) => EXP_out_1_port, 
                           EXP_out(0) => EXP_out_0_port);
   I3 : PackFP port map( SIGN => SIGN_out, EXP(7) => EXP_out_7_port, EXP(6) => 
                           EXP_out_6_port, EXP(5) => EXP_out_5_port, EXP(4) => 
                           EXP_out_4_port, EXP(3) => EXP_out_3_port, EXP(2) => 
                           EXP_out_2_port, EXP(1) => EXP_out_1_port, EXP(0) => 
                           EXP_out_0_port, SIG(22) => SIG_out_22_port, SIG(21) 
                           => SIG_out_21_port, SIG(20) => SIG_out_20_port, 
                           SIG(19) => SIG_out_19_port, SIG(18) => 
                           SIG_out_18_port, SIG(17) => SIG_out_17_port, SIG(16)
                           => SIG_out_16_port, SIG(15) => SIG_out_15_port, 
                           SIG(14) => SIG_out_14_port, SIG(13) => 
                           SIG_out_13_port, SIG(12) => SIG_out_12_port, SIG(11)
                           => SIG_out_11_port, SIG(10) => SIG_out_10_port, 
                           SIG(9) => SIG_out_9_port, SIG(8) => SIG_out_8_port, 
                           SIG(7) => SIG_out_7_port, SIG(6) => SIG_out_6_port, 
                           SIG(5) => SIG_out_5_port, SIG(4) => SIG_out_4_port, 
                           SIG(3) => SIG_out_3_port, SIG(2) => SIG_out_2_port, 
                           SIG(1) => SIG_out_1_port, SIG(0) => SIG_out_0_port, 
                           isNaN => isNaN, isINF => isINF, isZ => n33, FP(31) 
                           => FP_31_port, FP(30) => FP_30_port, FP(29) => 
                           FP_29_port, FP(28) => FP_28_port, FP(27) => 
                           FP_27_port, FP(26) => FP_26_port, FP(25) => 
                           FP_25_port, FP(24) => FP_24_port, FP(23) => 
                           FP_23_port, FP(22) => FP_22_port, FP(21) => 
                           FP_21_port, FP(20) => FP_20_port, FP(19) => 
                           FP_19_port, FP(18) => FP_18_port, FP(17) => 
                           FP_17_port, FP(16) => FP_16_port, FP(15) => 
                           FP_15_port, FP(14) => FP_14_port, FP(13) => 
                           FP_13_port, FP(12) => FP_12_port, FP(11) => 
                           FP_11_port, FP(10) => FP_10_port, FP(9) => FP_9_port
                           , FP(8) => FP_8_port, FP(7) => FP_7_port, FP(6) => 
                           FP_6_port, FP(5) => FP_5_port, FP(4) => FP_4_port, 
                           FP(3) => FP_3_port, FP(2) => FP_2_port, FP(1) => 
                           FP_1_port, FP(0) => FP_0_port);
   FP_Z_reg_31_inst : DFF_X1 port map( D => FP_31_port, CK => clk, Q => 
                           FP_Z(31), QN => n_1049);
   FP_Z_reg_30_inst : DFF_X1 port map( D => FP_30_port, CK => clk, Q => 
                           FP_Z(30), QN => n_1050);
   FP_Z_reg_29_inst : DFF_X1 port map( D => FP_29_port, CK => clk, Q => 
                           FP_Z(29), QN => n_1051);
   FP_Z_reg_28_inst : DFF_X1 port map( D => FP_28_port, CK => clk, Q => 
                           FP_Z(28), QN => n_1052);
   FP_Z_reg_27_inst : DFF_X1 port map( D => FP_27_port, CK => clk, Q => 
                           FP_Z(27), QN => n_1053);
   FP_Z_reg_26_inst : DFF_X1 port map( D => FP_26_port, CK => clk, Q => 
                           FP_Z(26), QN => n_1054);
   FP_Z_reg_25_inst : DFF_X1 port map( D => FP_25_port, CK => clk, Q => 
                           FP_Z(25), QN => n_1055);
   FP_Z_reg_24_inst : DFF_X1 port map( D => FP_24_port, CK => clk, Q => 
                           FP_Z(24), QN => n_1056);
   FP_Z_reg_23_inst : DFF_X1 port map( D => FP_23_port, CK => clk, Q => 
                           FP_Z(23), QN => n_1057);
   FP_Z_reg_22_inst : DFF_X1 port map( D => FP_22_port, CK => clk, Q => 
                           FP_Z(22), QN => n_1058);
   FP_Z_reg_21_inst : DFF_X1 port map( D => FP_21_port, CK => clk, Q => 
                           FP_Z(21), QN => n_1059);
   FP_Z_reg_20_inst : DFF_X1 port map( D => FP_20_port, CK => clk, Q => 
                           FP_Z(20), QN => n_1060);
   FP_Z_reg_19_inst : DFF_X1 port map( D => FP_19_port, CK => clk, Q => 
                           FP_Z(19), QN => n_1061);
   FP_Z_reg_18_inst : DFF_X1 port map( D => FP_18_port, CK => clk, Q => 
                           FP_Z(18), QN => n_1062);
   FP_Z_reg_17_inst : DFF_X1 port map( D => FP_17_port, CK => clk, Q => 
                           FP_Z(17), QN => n_1063);
   FP_Z_reg_16_inst : DFF_X1 port map( D => FP_16_port, CK => clk, Q => 
                           FP_Z(16), QN => n_1064);
   FP_Z_reg_15_inst : DFF_X1 port map( D => FP_15_port, CK => clk, Q => 
                           FP_Z(15), QN => n_1065);
   FP_Z_reg_14_inst : DFF_X1 port map( D => FP_14_port, CK => clk, Q => 
                           FP_Z(14), QN => n_1066);
   FP_Z_reg_13_inst : DFF_X1 port map( D => FP_13_port, CK => clk, Q => 
                           FP_Z(13), QN => n_1067);
   FP_Z_reg_12_inst : DFF_X1 port map( D => FP_12_port, CK => clk, Q => 
                           FP_Z(12), QN => n_1068);
   FP_Z_reg_11_inst : DFF_X1 port map( D => FP_11_port, CK => clk, Q => 
                           FP_Z(11), QN => n_1069);
   FP_Z_reg_10_inst : DFF_X1 port map( D => FP_10_port, CK => clk, Q => 
                           FP_Z(10), QN => n_1070);
   FP_Z_reg_9_inst : DFF_X1 port map( D => FP_9_port, CK => clk, Q => FP_Z(9), 
                           QN => n_1071);
   FP_Z_reg_8_inst : DFF_X1 port map( D => FP_8_port, CK => clk, Q => FP_Z(8), 
                           QN => n_1072);
   FP_Z_reg_7_inst : DFF_X1 port map( D => FP_7_port, CK => clk, Q => FP_Z(7), 
                           QN => n_1073);
   FP_Z_reg_6_inst : DFF_X1 port map( D => FP_6_port, CK => clk, Q => FP_Z(6), 
                           QN => n_1074);
   FP_Z_reg_5_inst : DFF_X1 port map( D => FP_5_port, CK => clk, Q => FP_Z(5), 
                           QN => n_1075);
   FP_Z_reg_4_inst : DFF_X1 port map( D => FP_4_port, CK => clk, Q => FP_Z(4), 
                           QN => n_1076);
   FP_Z_reg_3_inst : DFF_X1 port map( D => FP_3_port, CK => clk, Q => FP_Z(3), 
                           QN => n_1077);
   FP_Z_reg_2_inst : DFF_X1 port map( D => FP_2_port, CK => clk, Q => FP_Z(2), 
                           QN => n_1078);
   FP_Z_reg_1_inst : DFF_X1 port map( D => FP_1_port, CK => clk, Q => FP_Z(1), 
                           QN => n_1079);
   FP_Z_reg_0_inst : DFF_X1 port map( D => FP_0_port, CK => clk, Q => FP_Z(0), 
                           QN => n_1080);
   U3 : NOR2_X1 port map( A1 => n23, A2 => n22, ZN => n27);
   U4 : NAND2_X1 port map( A1 => EXP_out_3_port, A2 => EXP_out_4_port, ZN => 
                           n23);
   U5 : NAND2_X1 port map( A1 => EXP_out_5_port, A2 => EXP_out_6_port, ZN => 
                           n22);
   U6 : INV_X1 port map( A => EXP_out_0_port, ZN => n24);
   U7 : INV_X1 port map( A => EXP_out_2_port, ZN => n25);
   U8 : AOI21_X1 port map( B1 => n32, B2 => n31, A => n33, ZN => isINF);
   U9 : INV_X1 port map( A => isINF_tab, ZN => n31);
   U10 : INV_X1 port map( A => EXP_pos, ZN => n29);
   U11 : NOR2_X1 port map( A1 => n25, A2 => n24, ZN => n26);
   U12 : INV_X1 port map( A => SIG_out_5_port, ZN => n4);
   U13 : INV_X1 port map( A => SIG_out_4_port, ZN => n3);
   U14 : INV_X1 port map( A => SIG_out_3_port, ZN => n2);
   U15 : NOR3_X1 port map( A1 => SIG_out_0_port, A2 => SIG_out_1_port, A3 => 
                           SIG_out_2_port, ZN => n1);
   U16 : NAND4_X1 port map( A1 => n4, A2 => n3, A3 => n2, A4 => n1, ZN => n20);
   U17 : INV_X1 port map( A => SIG_out_11_port, ZN => n8);
   U18 : INV_X1 port map( A => SIG_out_10_port, ZN => n7);
   U19 : INV_X1 port map( A => SIG_out_9_port, ZN => n6);
   U20 : NOR3_X1 port map( A1 => SIG_out_6_port, A2 => SIG_out_7_port, A3 => 
                           SIG_out_8_port, ZN => n5);
   U21 : NAND4_X1 port map( A1 => n8, A2 => n7, A3 => n6, A4 => n5, ZN => n19);
   U22 : INV_X1 port map( A => SIG_out_17_port, ZN => n12);
   U23 : INV_X1 port map( A => SIG_out_16_port, ZN => n11);
   U24 : INV_X1 port map( A => SIG_out_15_port, ZN => n10);
   U25 : NOR3_X1 port map( A1 => SIG_out_12_port, A2 => SIG_out_13_port, A3 => 
                           SIG_out_14_port, ZN => n9);
   U26 : NAND4_X1 port map( A1 => n12, A2 => n11, A3 => n10, A4 => n9, ZN => 
                           n18);
   U27 : INV_X1 port map( A => SIG_out_20_port, ZN => n16);
   U28 : INV_X1 port map( A => SIG_out_19_port, ZN => n15);
   U29 : INV_X1 port map( A => SIG_out_18_port, ZN => n14);
   U30 : NOR3_X1 port map( A1 => SIG_out_21_port, A2 => SIG_out_22_port, A3 => 
                           SIG_out_norm2_26_port, ZN => n13);
   U31 : NAND4_X1 port map( A1 => n16, A2 => n15, A3 => n14, A4 => n13, ZN => 
                           n17);
   U32 : NOR4_X1 port map( A1 => n20, A2 => n19, A3 => n18, A4 => n17, ZN => 
                           n21);
   U33 : AOI211_X1 port map( C1 => EXP_out_7_port, C2 => EXP_neg, A => isZ_tab,
                           B => n21, ZN => n30);
   U34 : INV_X1 port map( A => n30, ZN => n33);
   U35 : NAND3_X1 port map( A1 => EXP_out_1_port, A2 => n27, A3 => n26, ZN => 
                           n28);
   U36 : MUX2_X1 port map( A => n29, B => n28, S => EXP_out_7_port, Z => n32);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage3 is

   port( EXP_in : in std_logic_vector (7 downto 0);  EXP_neg_stage2, 
         EXP_pos_stage2, SIGN_out_stage2 : in std_logic;  SIG_in : in 
         std_logic_vector (27 downto 0);  clk, isINF_stage2, isNaN_stage2, 
         isZ_tab_stage2 : in std_logic;  EXP_neg : out std_logic;  
         EXP_out_round : out std_logic_vector (7 downto 0);  EXP_pos, SIGN_out 
         : out std_logic;  SIG_out_round : out std_logic_vector (27 downto 0); 
         isINF_tab, isNaN, isZ_tab : out std_logic);

end FPmul_stage3;

architecture SYN_struct of FPmul_stage3 is

   component FPround_SIG_width28
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0));
   end component;
   
   component FPnormalize_SIG_width28_0
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0));
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal EXP_out_7_port, EXP_out_6_port, EXP_out_5_port, EXP_out_4_port, 
      EXP_out_3_port, EXP_out_2_port, EXP_out_1_port, EXP_out_0_port, 
      SIG_out_27_port, SIG_out_26_port, SIG_out_25_port, SIG_out_24_port, 
      SIG_out_23_port, SIG_out_22_port, SIG_out_21_port, SIG_out_20_port, 
      SIG_out_19_port, SIG_out_18_port, SIG_out_17_port, SIG_out_16_port, 
      SIG_out_15_port, SIG_out_14_port, SIG_out_13_port, SIG_out_12_port, 
      SIG_out_11_port, SIG_out_10_port, SIG_out_9_port, SIG_out_8_port, 
      SIG_out_7_port, SIG_out_6_port, SIG_out_5_port, SIG_out_4_port, 
      SIG_out_3_port, SIG_out_1_port, SIG_out_0_port, SIG_out_norm_27_port, 
      SIG_out_norm_26_port, SIG_out_norm_25_port, SIG_out_norm_24_port, 
      SIG_out_norm_23_port, SIG_out_norm_22_port, SIG_out_norm_21_port, 
      SIG_out_norm_20_port, SIG_out_norm_19_port, SIG_out_norm_18_port, 
      SIG_out_norm_17_port, SIG_out_norm_16_port, SIG_out_norm_15_port, 
      SIG_out_norm_14_port, SIG_out_norm_13_port, SIG_out_norm_12_port, 
      SIG_out_norm_11_port, SIG_out_norm_10_port, SIG_out_norm_9_port, 
      SIG_out_norm_8_port, SIG_out_norm_7_port, SIG_out_norm_6_port, 
      SIG_out_norm_5_port, SIG_out_norm_4_port, SIG_out_norm_3_port, 
      SIG_out_norm_2_port, SIG_out_norm_1_port, SIG_out_norm_0_port, 
      EXP_out_norm_7_port, EXP_out_norm_6_port, EXP_out_norm_5_port, 
      EXP_out_norm_4_port, EXP_out_norm_3_port, EXP_out_norm_2_port, 
      EXP_out_norm_1_port, EXP_out_norm_0_port, n_1081, n_1082, n_1083, n_1084,
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123 : std_logic;

begin
   
   EXP_out_round_reg_7_inst : DFF_X1 port map( D => EXP_out_7_port, CK => clk, 
                           Q => EXP_out_round(7), QN => n_1081);
   EXP_out_round_reg_6_inst : DFF_X1 port map( D => EXP_out_6_port, CK => clk, 
                           Q => EXP_out_round(6), QN => n_1082);
   EXP_out_round_reg_5_inst : DFF_X1 port map( D => EXP_out_5_port, CK => clk, 
                           Q => EXP_out_round(5), QN => n_1083);
   EXP_out_round_reg_4_inst : DFF_X1 port map( D => EXP_out_4_port, CK => clk, 
                           Q => EXP_out_round(4), QN => n_1084);
   EXP_out_round_reg_3_inst : DFF_X1 port map( D => EXP_out_3_port, CK => clk, 
                           Q => EXP_out_round(3), QN => n_1085);
   EXP_out_round_reg_2_inst : DFF_X1 port map( D => EXP_out_2_port, CK => clk, 
                           Q => EXP_out_round(2), QN => n_1086);
   EXP_out_round_reg_1_inst : DFF_X1 port map( D => EXP_out_1_port, CK => clk, 
                           Q => EXP_out_round(1), QN => n_1087);
   EXP_out_round_reg_0_inst : DFF_X1 port map( D => EXP_out_0_port, CK => clk, 
                           Q => EXP_out_round(0), QN => n_1088);
   SIG_out_round_reg_27_inst : DFF_X1 port map( D => SIG_out_27_port, CK => clk
                           , Q => SIG_out_round(27), QN => n_1089);
   SIG_out_round_reg_26_inst : DFF_X1 port map( D => SIG_out_26_port, CK => clk
                           , Q => SIG_out_round(26), QN => n_1090);
   SIG_out_round_reg_25_inst : DFF_X1 port map( D => SIG_out_25_port, CK => clk
                           , Q => SIG_out_round(25), QN => n_1091);
   SIG_out_round_reg_24_inst : DFF_X1 port map( D => SIG_out_24_port, CK => clk
                           , Q => SIG_out_round(24), QN => n_1092);
   SIG_out_round_reg_23_inst : DFF_X1 port map( D => SIG_out_23_port, CK => clk
                           , Q => SIG_out_round(23), QN => n_1093);
   SIG_out_round_reg_22_inst : DFF_X1 port map( D => SIG_out_22_port, CK => clk
                           , Q => SIG_out_round(22), QN => n_1094);
   SIG_out_round_reg_21_inst : DFF_X1 port map( D => SIG_out_21_port, CK => clk
                           , Q => SIG_out_round(21), QN => n_1095);
   SIG_out_round_reg_20_inst : DFF_X1 port map( D => SIG_out_20_port, CK => clk
                           , Q => SIG_out_round(20), QN => n_1096);
   SIG_out_round_reg_19_inst : DFF_X1 port map( D => SIG_out_19_port, CK => clk
                           , Q => SIG_out_round(19), QN => n_1097);
   SIG_out_round_reg_18_inst : DFF_X1 port map( D => SIG_out_18_port, CK => clk
                           , Q => SIG_out_round(18), QN => n_1098);
   SIG_out_round_reg_17_inst : DFF_X1 port map( D => SIG_out_17_port, CK => clk
                           , Q => SIG_out_round(17), QN => n_1099);
   SIG_out_round_reg_16_inst : DFF_X1 port map( D => SIG_out_16_port, CK => clk
                           , Q => SIG_out_round(16), QN => n_1100);
   SIG_out_round_reg_15_inst : DFF_X1 port map( D => SIG_out_15_port, CK => clk
                           , Q => SIG_out_round(15), QN => n_1101);
   SIG_out_round_reg_14_inst : DFF_X1 port map( D => SIG_out_14_port, CK => clk
                           , Q => SIG_out_round(14), QN => n_1102);
   SIG_out_round_reg_13_inst : DFF_X1 port map( D => SIG_out_13_port, CK => clk
                           , Q => SIG_out_round(13), QN => n_1103);
   SIG_out_round_reg_12_inst : DFF_X1 port map( D => SIG_out_12_port, CK => clk
                           , Q => SIG_out_round(12), QN => n_1104);
   SIG_out_round_reg_11_inst : DFF_X1 port map( D => SIG_out_11_port, CK => clk
                           , Q => SIG_out_round(11), QN => n_1105);
   SIG_out_round_reg_10_inst : DFF_X1 port map( D => SIG_out_10_port, CK => clk
                           , Q => SIG_out_round(10), QN => n_1106);
   SIG_out_round_reg_9_inst : DFF_X1 port map( D => SIG_out_9_port, CK => clk, 
                           Q => SIG_out_round(9), QN => n_1107);
   SIG_out_round_reg_8_inst : DFF_X1 port map( D => SIG_out_8_port, CK => clk, 
                           Q => SIG_out_round(8), QN => n_1108);
   SIG_out_round_reg_7_inst : DFF_X1 port map( D => SIG_out_7_port, CK => clk, 
                           Q => SIG_out_round(7), QN => n_1109);
   SIG_out_round_reg_6_inst : DFF_X1 port map( D => SIG_out_6_port, CK => clk, 
                           Q => SIG_out_round(6), QN => n_1110);
   SIG_out_round_reg_5_inst : DFF_X1 port map( D => SIG_out_5_port, CK => clk, 
                           Q => SIG_out_round(5), QN => n_1111);
   SIG_out_round_reg_4_inst : DFF_X1 port map( D => SIG_out_4_port, CK => clk, 
                           Q => SIG_out_round(4), QN => n_1112);
   SIG_out_round_reg_3_inst : DFF_X1 port map( D => SIG_out_3_port, CK => clk, 
                           Q => SIG_out_round(3), QN => n_1113);
   SIG_out_round_reg_1_inst : DFF_X1 port map( D => SIG_out_1_port, CK => clk, 
                           Q => SIG_out_round(1), QN => n_1114);
   SIG_out_round_reg_0_inst : DFF_X1 port map( D => SIG_out_0_port, CK => clk, 
                           Q => SIG_out_round(0), QN => n_1115);
   isINF_tab_reg : DFF_X1 port map( D => isINF_stage2, CK => clk, Q => 
                           isINF_tab, QN => n_1116);
   isNaN_reg : DFF_X1 port map( D => isNaN_stage2, CK => clk, Q => isNaN, QN =>
                           n_1117);
   isZ_tab_reg : DFF_X1 port map( D => isZ_tab_stage2, CK => clk, Q => isZ_tab,
                           QN => n_1118);
   SIGN_out_reg : DFF_X1 port map( D => SIGN_out_stage2, CK => clk, Q => 
                           SIGN_out, QN => n_1119);
   EXP_pos_reg : DFF_X1 port map( D => EXP_pos_stage2, CK => clk, Q => EXP_pos,
                           QN => n_1120);
   EXP_neg_reg : DFF_X1 port map( D => EXP_neg_stage2, CK => clk, Q => EXP_neg,
                           QN => n_1121);
   I9 : FPnormalize_SIG_width28_0 port map( SIG_in(27) => SIG_in(27), 
                           SIG_in(26) => SIG_in(26), SIG_in(25) => SIG_in(25), 
                           SIG_in(24) => SIG_in(24), SIG_in(23) => SIG_in(23), 
                           SIG_in(22) => SIG_in(22), SIG_in(21) => SIG_in(21), 
                           SIG_in(20) => SIG_in(20), SIG_in(19) => SIG_in(19), 
                           SIG_in(18) => SIG_in(18), SIG_in(17) => SIG_in(17), 
                           SIG_in(16) => SIG_in(16), SIG_in(15) => SIG_in(15), 
                           SIG_in(14) => SIG_in(14), SIG_in(13) => SIG_in(13), 
                           SIG_in(12) => SIG_in(12), SIG_in(11) => SIG_in(11), 
                           SIG_in(10) => SIG_in(10), SIG_in(9) => SIG_in(9), 
                           SIG_in(8) => SIG_in(8), SIG_in(7) => SIG_in(7), 
                           SIG_in(6) => SIG_in(6), SIG_in(5) => SIG_in(5), 
                           SIG_in(4) => SIG_in(4), SIG_in(3) => SIG_in(3), 
                           SIG_in(2) => SIG_in(2), SIG_in(1) => SIG_in(1), 
                           SIG_in(0) => SIG_in(0), EXP_in(7) => EXP_in(7), 
                           EXP_in(6) => EXP_in(6), EXP_in(5) => EXP_in(5), 
                           EXP_in(4) => EXP_in(4), EXP_in(3) => EXP_in(3), 
                           EXP_in(2) => EXP_in(2), EXP_in(1) => EXP_in(1), 
                           EXP_in(0) => EXP_in(0), SIG_out(27) => n_1122, 
                           SIG_out(26) => SIG_out_norm_26_port, SIG_out(25) => 
                           SIG_out_norm_25_port, SIG_out(24) => 
                           SIG_out_norm_24_port, SIG_out(23) => 
                           SIG_out_norm_23_port, SIG_out(22) => 
                           SIG_out_norm_22_port, SIG_out(21) => 
                           SIG_out_norm_21_port, SIG_out(20) => 
                           SIG_out_norm_20_port, SIG_out(19) => 
                           SIG_out_norm_19_port, SIG_out(18) => 
                           SIG_out_norm_18_port, SIG_out(17) => 
                           SIG_out_norm_17_port, SIG_out(16) => 
                           SIG_out_norm_16_port, SIG_out(15) => 
                           SIG_out_norm_15_port, SIG_out(14) => 
                           SIG_out_norm_14_port, SIG_out(13) => 
                           SIG_out_norm_13_port, SIG_out(12) => 
                           SIG_out_norm_12_port, SIG_out(11) => 
                           SIG_out_norm_11_port, SIG_out(10) => 
                           SIG_out_norm_10_port, SIG_out(9) => 
                           SIG_out_norm_9_port, SIG_out(8) => 
                           SIG_out_norm_8_port, SIG_out(7) => 
                           SIG_out_norm_7_port, SIG_out(6) => 
                           SIG_out_norm_6_port, SIG_out(5) => 
                           SIG_out_norm_5_port, SIG_out(4) => 
                           SIG_out_norm_4_port, SIG_out(3) => 
                           SIG_out_norm_3_port, SIG_out(2) => 
                           SIG_out_norm_2_port, SIG_out(1) => 
                           SIG_out_norm_1_port, SIG_out(0) => 
                           SIG_out_norm_0_port, EXP_out(7) => 
                           EXP_out_norm_7_port, EXP_out(6) => 
                           EXP_out_norm_6_port, EXP_out(5) => 
                           EXP_out_norm_5_port, EXP_out(4) => 
                           EXP_out_norm_4_port, EXP_out(3) => 
                           EXP_out_norm_3_port, EXP_out(2) => 
                           EXP_out_norm_2_port, EXP_out(1) => 
                           EXP_out_norm_1_port, EXP_out(0) => 
                           EXP_out_norm_0_port);
   I11 : FPround_SIG_width28 port map( SIG_in(27) => SIG_out_norm_27_port, 
                           SIG_in(26) => SIG_out_norm_26_port, SIG_in(25) => 
                           SIG_out_norm_25_port, SIG_in(24) => 
                           SIG_out_norm_24_port, SIG_in(23) => 
                           SIG_out_norm_23_port, SIG_in(22) => 
                           SIG_out_norm_22_port, SIG_in(21) => 
                           SIG_out_norm_21_port, SIG_in(20) => 
                           SIG_out_norm_20_port, SIG_in(19) => 
                           SIG_out_norm_19_port, SIG_in(18) => 
                           SIG_out_norm_18_port, SIG_in(17) => 
                           SIG_out_norm_17_port, SIG_in(16) => 
                           SIG_out_norm_16_port, SIG_in(15) => 
                           SIG_out_norm_15_port, SIG_in(14) => 
                           SIG_out_norm_14_port, SIG_in(13) => 
                           SIG_out_norm_13_port, SIG_in(12) => 
                           SIG_out_norm_12_port, SIG_in(11) => 
                           SIG_out_norm_11_port, SIG_in(10) => 
                           SIG_out_norm_10_port, SIG_in(9) => 
                           SIG_out_norm_9_port, SIG_in(8) => 
                           SIG_out_norm_8_port, SIG_in(7) => 
                           SIG_out_norm_7_port, SIG_in(6) => 
                           SIG_out_norm_6_port, SIG_in(5) => 
                           SIG_out_norm_5_port, SIG_in(4) => 
                           SIG_out_norm_4_port, SIG_in(3) => 
                           SIG_out_norm_3_port, SIG_in(2) => 
                           SIG_out_norm_2_port, SIG_in(1) => 
                           SIG_out_norm_1_port, SIG_in(0) => 
                           SIG_out_norm_0_port, EXP_in(7) => 
                           EXP_out_norm_7_port, EXP_in(6) => 
                           EXP_out_norm_6_port, EXP_in(5) => 
                           EXP_out_norm_5_port, EXP_in(4) => 
                           EXP_out_norm_4_port, EXP_in(3) => 
                           EXP_out_norm_3_port, EXP_in(2) => 
                           EXP_out_norm_2_port, EXP_in(1) => 
                           EXP_out_norm_1_port, EXP_in(0) => 
                           EXP_out_norm_0_port, SIG_out(27) => SIG_out_27_port,
                           SIG_out(26) => SIG_out_26_port, SIG_out(25) => 
                           SIG_out_25_port, SIG_out(24) => SIG_out_24_port, 
                           SIG_out(23) => SIG_out_23_port, SIG_out(22) => 
                           SIG_out_22_port, SIG_out(21) => SIG_out_21_port, 
                           SIG_out(20) => SIG_out_20_port, SIG_out(19) => 
                           SIG_out_19_port, SIG_out(18) => SIG_out_18_port, 
                           SIG_out(17) => SIG_out_17_port, SIG_out(16) => 
                           SIG_out_16_port, SIG_out(15) => SIG_out_15_port, 
                           SIG_out(14) => SIG_out_14_port, SIG_out(13) => 
                           SIG_out_13_port, SIG_out(12) => SIG_out_12_port, 
                           SIG_out(11) => SIG_out_11_port, SIG_out(10) => 
                           SIG_out_10_port, SIG_out(9) => SIG_out_9_port, 
                           SIG_out(8) => SIG_out_8_port, SIG_out(7) => 
                           SIG_out_7_port, SIG_out(6) => SIG_out_6_port, 
                           SIG_out(5) => SIG_out_5_port, SIG_out(4) => 
                           SIG_out_4_port, SIG_out(3) => SIG_out_3_port, 
                           SIG_out(2) => n_1123, SIG_out(1) => SIG_out_1_port, 
                           SIG_out(0) => SIG_out_0_port, EXP_out(7) => 
                           EXP_out_7_port, EXP_out(6) => EXP_out_6_port, 
                           EXP_out(5) => EXP_out_5_port, EXP_out(4) => 
                           EXP_out_4_port, EXP_out(3) => EXP_out_3_port, 
                           EXP_out(2) => EXP_out_2_port, EXP_out(1) => 
                           EXP_out_1_port, EXP_out(0) => EXP_out_0_port);
   SIG_out_round(2) <= '0';
   SIG_out_norm_27_port <= '0';

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage2 is

   port( A_EXP : in std_logic_vector (7 downto 0);  A_SIG : in std_logic_vector
         (31 downto 0);  B_EXP : in std_logic_vector (7 downto 0);  B_SIG : in 
         std_logic_vector (31 downto 0);  SIGN_out_stage1, clk, isINF_stage1, 
         isNaN_stage1, isZ_tab_stage1 : in std_logic;  EXP_in : out 
         std_logic_vector (7 downto 0);  EXP_neg_stage2, EXP_pos_stage2, 
         SIGN_out_stage2 : out std_logic;  SIG_in : out std_logic_vector (27 
         downto 0);  isINF_stage2, isNaN_stage2, isZ_tab_stage2 : out std_logic
         );

end FPmul_stage2;

architecture SYN_struct of FPmul_stage2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FPmul_stage2_DW01_add_0
      port( A, B : in std_logic_vector (7 downto 0);  CI : in std_logic;  SUM :
            out std_logic_vector (7 downto 0);  CO : out std_logic);
   end component;
   
   component MBE
      port( A, B : in std_logic_vector (31 downto 0);  C : out std_logic_vector
            (63 downto 0));
   end component;
   
   signal X_Logic1_port, SIG_in_int_27_port, SIG_in_int_26_port, 
      SIG_in_int_25_port, SIG_in_int_24_port, SIG_in_int_23_port, 
      SIG_in_int_22_port, SIG_in_int_21_port, SIG_in_int_20_port, 
      SIG_in_int_19_port, SIG_in_int_18_port, SIG_in_int_17_port, 
      SIG_in_int_16_port, SIG_in_int_15_port, SIG_in_int_14_port, 
      SIG_in_int_13_port, SIG_in_int_12_port, SIG_in_int_11_port, 
      SIG_in_int_10_port, SIG_in_int_9_port, SIG_in_int_8_port, 
      SIG_in_int_7_port, SIG_in_int_6_port, SIG_in_int_5_port, 
      SIG_in_int_4_port, SIG_in_int_3_port, SIG_in_int_2_port, 
      SIG_in_int_1_port, SIG_in_int_0_port, EXP_pos_int, N0, mw_I4sum_7_port, 
      mw_I4sum_6_port, mw_I4sum_5_port, mw_I4sum_4_port, mw_I4sum_3_port, 
      mw_I4sum_2_port, mw_I4sum_1_port, mw_I4sum_0_port, n1, n2, n3, n4, n5, n6
      , n7, n8, n9, n10, n11, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202 : std_logic;

begin
   
   X_Logic1_port <= '1';
   EXP_in_reg_7_inst : DFF_X1 port map( D => n11, CK => clk, Q => EXP_in(7), QN
                           => n_1124);
   EXP_in_reg_6_inst : DFF_X1 port map( D => mw_I4sum_6_port, CK => clk, Q => 
                           EXP_in(6), QN => n_1125);
   EXP_in_reg_5_inst : DFF_X1 port map( D => mw_I4sum_5_port, CK => clk, Q => 
                           EXP_in(5), QN => n_1126);
   EXP_in_reg_4_inst : DFF_X1 port map( D => mw_I4sum_4_port, CK => clk, Q => 
                           EXP_in(4), QN => n_1127);
   EXP_in_reg_3_inst : DFF_X1 port map( D => mw_I4sum_3_port, CK => clk, Q => 
                           EXP_in(3), QN => n_1128);
   EXP_in_reg_2_inst : DFF_X1 port map( D => mw_I4sum_2_port, CK => clk, Q => 
                           EXP_in(2), QN => n_1129);
   EXP_in_reg_1_inst : DFF_X1 port map( D => mw_I4sum_1_port, CK => clk, Q => 
                           EXP_in(1), QN => n_1130);
   EXP_in_reg_0_inst : DFF_X1 port map( D => mw_I4sum_0_port, CK => clk, Q => 
                           EXP_in(0), QN => n_1131);
   EXP_pos_stage2_reg : DFF_X1 port map( D => EXP_pos_int, CK => clk, Q => 
                           EXP_pos_stage2, QN => n_1132);
   EXP_neg_stage2_reg : DFF_X1 port map( D => N0, CK => clk, Q => 
                           EXP_neg_stage2, QN => n_1133);
   isINF_stage2_reg : DFF_X1 port map( D => isINF_stage1, CK => clk, Q => 
                           isINF_stage2, QN => n_1134);
   isNaN_stage2_reg : DFF_X1 port map( D => isNaN_stage1, CK => clk, Q => 
                           isNaN_stage2, QN => n_1135);
   isZ_tab_stage2_reg : DFF_X1 port map( D => isZ_tab_stage1, CK => clk, Q => 
                           isZ_tab_stage2, QN => n_1136);
   SIGN_out_stage2_reg : DFF_X1 port map( D => SIGN_out_stage1, CK => clk, Q =>
                           SIGN_out_stage2, QN => n_1137);
   MBE_SIG : MBE port map( A(31) => A_SIG(31), A(30) => A_SIG(30), A(29) => 
                           A_SIG(29), A(28) => A_SIG(28), A(27) => A_SIG(27), 
                           A(26) => A_SIG(26), A(25) => A_SIG(25), A(24) => 
                           A_SIG(24), A(23) => A_SIG(23), A(22) => A_SIG(22), 
                           A(21) => A_SIG(21), A(20) => A_SIG(20), A(19) => 
                           A_SIG(19), A(18) => A_SIG(18), A(17) => A_SIG(17), 
                           A(16) => A_SIG(16), A(15) => A_SIG(15), A(14) => 
                           A_SIG(14), A(13) => A_SIG(13), A(12) => A_SIG(12), 
                           A(11) => A_SIG(11), A(10) => A_SIG(10), A(9) => 
                           A_SIG(9), A(8) => A_SIG(8), A(7) => A_SIG(7), A(6) 
                           => A_SIG(6), A(5) => A_SIG(5), A(4) => A_SIG(4), 
                           A(3) => A_SIG(3), A(2) => A_SIG(2), A(1) => A_SIG(1)
                           , A(0) => A_SIG(0), B(31) => B_SIG(31), B(30) => 
                           B_SIG(30), B(29) => B_SIG(29), B(28) => B_SIG(28), 
                           B(27) => B_SIG(27), B(26) => B_SIG(26), B(25) => 
                           B_SIG(25), B(24) => B_SIG(24), B(23) => B_SIG(23), 
                           B(22) => B_SIG(22), B(21) => B_SIG(21), B(20) => 
                           B_SIG(20), B(19) => B_SIG(19), B(18) => B_SIG(18), 
                           B(17) => B_SIG(17), B(16) => B_SIG(16), B(15) => 
                           B_SIG(15), B(14) => B_SIG(14), B(13) => B_SIG(13), 
                           B(12) => B_SIG(12), B(11) => B_SIG(11), B(10) => 
                           B_SIG(10), B(9) => B_SIG(9), B(8) => B_SIG(8), B(7) 
                           => B_SIG(7), B(6) => B_SIG(6), B(5) => B_SIG(5), 
                           B(4) => B_SIG(4), B(3) => B_SIG(3), B(2) => B_SIG(2)
                           , B(1) => B_SIG(1), B(0) => B_SIG(0), C(63) => 
                           n_1138, C(62) => n_1139, C(61) => n_1140, C(60) => 
                           n_1141, C(59) => n_1142, C(58) => n_1143, C(57) => 
                           n_1144, C(56) => n_1145, C(55) => n_1146, C(54) => 
                           n_1147, C(53) => n_1148, C(52) => n_1149, C(51) => 
                           n_1150, C(50) => n_1151, C(49) => n_1152, C(48) => 
                           n_1153, C(47) => SIG_in_int_27_port, C(46) => 
                           SIG_in_int_26_port, C(45) => SIG_in_int_25_port, 
                           C(44) => SIG_in_int_24_port, C(43) => 
                           SIG_in_int_23_port, C(42) => SIG_in_int_22_port, 
                           C(41) => SIG_in_int_21_port, C(40) => 
                           SIG_in_int_20_port, C(39) => SIG_in_int_19_port, 
                           C(38) => SIG_in_int_18_port, C(37) => 
                           SIG_in_int_17_port, C(36) => SIG_in_int_16_port, 
                           C(35) => SIG_in_int_15_port, C(34) => 
                           SIG_in_int_14_port, C(33) => SIG_in_int_13_port, 
                           C(32) => SIG_in_int_12_port, C(31) => 
                           SIG_in_int_11_port, C(30) => SIG_in_int_10_port, 
                           C(29) => SIG_in_int_9_port, C(28) => 
                           SIG_in_int_8_port, C(27) => SIG_in_int_7_port, C(26)
                           => SIG_in_int_6_port, C(25) => SIG_in_int_5_port, 
                           C(24) => SIG_in_int_4_port, C(23) => 
                           SIG_in_int_3_port, C(22) => SIG_in_int_2_port, C(21)
                           => SIG_in_int_1_port, C(20) => SIG_in_int_0_port, 
                           C(19) => n_1154, C(18) => n_1155, C(17) => n_1156, 
                           C(16) => n_1157, C(15) => n_1158, C(14) => n_1159, 
                           C(13) => n_1160, C(12) => n_1161, C(11) => n_1162, 
                           C(10) => n_1163, C(9) => n_1164, C(8) => n_1165, 
                           C(7) => n_1166, C(6) => n_1167, C(5) => n_1168, C(4)
                           => n_1169, C(3) => n_1170, C(2) => n_1171, C(1) => 
                           n_1172, C(0) => n_1173);
   add_1_root_add_131_2 : FPmul_stage2_DW01_add_0 port map( A(7) => A_EXP(7), 
                           A(6) => A_EXP(6), A(5) => A_EXP(5), A(4) => A_EXP(4)
                           , A(3) => A_EXP(3), A(2) => A_EXP(2), A(1) => 
                           A_EXP(1), A(0) => A_EXP(0), B(7) => B_EXP(7), B(6) 
                           => B_EXP(6), B(5) => B_EXP(5), B(4) => B_EXP(4), 
                           B(3) => B_EXP(3), B(2) => B_EXP(2), B(1) => B_EXP(1)
                           , B(0) => B_EXP(0), CI => X_Logic1_port, SUM(7) => 
                           mw_I4sum_7_port, SUM(6) => mw_I4sum_6_port, SUM(5) 
                           => mw_I4sum_5_port, SUM(4) => mw_I4sum_4_port, 
                           SUM(3) => mw_I4sum_3_port, SUM(2) => mw_I4sum_2_port
                           , SUM(1) => mw_I4sum_1_port, SUM(0) => 
                           mw_I4sum_0_port, CO => n_1174);
   SIG_in_reg_11_inst : DFF_X1 port map( D => SIG_in_int_11_port, CK => clk, Q 
                           => SIG_in(11), QN => n_1175);
   SIG_in_reg_10_inst : DFF_X1 port map( D => SIG_in_int_10_port, CK => clk, Q 
                           => SIG_in(10), QN => n_1176);
   SIG_in_reg_9_inst : DFF_X1 port map( D => SIG_in_int_9_port, CK => clk, Q =>
                           SIG_in(9), QN => n_1177);
   SIG_in_reg_8_inst : DFF_X1 port map( D => SIG_in_int_8_port, CK => clk, Q =>
                           SIG_in(8), QN => n_1178);
   SIG_in_reg_3_inst : DFF_X1 port map( D => SIG_in_int_3_port, CK => clk, Q =>
                           SIG_in(3), QN => n_1179);
   SIG_in_reg_2_inst : DFF_X1 port map( D => SIG_in_int_2_port, CK => clk, Q =>
                           SIG_in(2), QN => n_1180);
   SIG_in_reg_1_inst : DFF_X1 port map( D => SIG_in_int_1_port, CK => clk, Q =>
                           SIG_in(1), QN => n_1181);
   SIG_in_reg_0_inst : DFF_X1 port map( D => SIG_in_int_0_port, CK => clk, Q =>
                           SIG_in(0), QN => n_1182);
   SIG_in_reg_7_inst : DFF_X1 port map( D => SIG_in_int_7_port, CK => clk, Q =>
                           SIG_in(7), QN => n_1183);
   SIG_in_reg_6_inst : DFF_X1 port map( D => SIG_in_int_6_port, CK => clk, Q =>
                           SIG_in(6), QN => n_1184);
   SIG_in_reg_5_inst : DFF_X1 port map( D => SIG_in_int_5_port, CK => clk, Q =>
                           SIG_in(5), QN => n_1185);
   SIG_in_reg_4_inst : DFF_X1 port map( D => SIG_in_int_4_port, CK => clk, Q =>
                           SIG_in(4), QN => n_1186);
   SIG_in_reg_14_inst : DFF_X1 port map( D => SIG_in_int_14_port, CK => clk, Q 
                           => SIG_in(14), QN => n_1187);
   SIG_in_reg_13_inst : DFF_X1 port map( D => SIG_in_int_13_port, CK => clk, Q 
                           => SIG_in(13), QN => n_1188);
   SIG_in_reg_12_inst : DFF_X1 port map( D => SIG_in_int_12_port, CK => clk, Q 
                           => SIG_in(12), QN => n_1189);
   SIG_in_reg_15_inst : DFF_X1 port map( D => SIG_in_int_15_port, CK => clk, Q 
                           => SIG_in(15), QN => n_1190);
   SIG_in_reg_26_inst : DFF_X1 port map( D => SIG_in_int_26_port, CK => clk, Q 
                           => SIG_in(26), QN => n_1191);
   SIG_in_reg_25_inst : DFF_X1 port map( D => SIG_in_int_25_port, CK => clk, Q 
                           => SIG_in(25), QN => n_1192);
   SIG_in_reg_24_inst : DFF_X1 port map( D => SIG_in_int_24_port, CK => clk, Q 
                           => SIG_in(24), QN => n_1193);
   SIG_in_reg_22_inst : DFF_X1 port map( D => SIG_in_int_22_port, CK => clk, Q 
                           => SIG_in(22), QN => n_1194);
   SIG_in_reg_21_inst : DFF_X1 port map( D => SIG_in_int_21_port, CK => clk, Q 
                           => SIG_in(21), QN => n_1195);
   SIG_in_reg_20_inst : DFF_X1 port map( D => SIG_in_int_20_port, CK => clk, Q 
                           => SIG_in(20), QN => n_1196);
   SIG_in_reg_18_inst : DFF_X1 port map( D => SIG_in_int_18_port, CK => clk, Q 
                           => SIG_in(18), QN => n_1197);
   SIG_in_reg_17_inst : DFF_X1 port map( D => SIG_in_int_17_port, CK => clk, Q 
                           => SIG_in(17), QN => n_1198);
   SIG_in_reg_16_inst : DFF_X1 port map( D => SIG_in_int_16_port, CK => clk, Q 
                           => SIG_in(16), QN => n_1199);
   SIG_in_reg_23_inst : DFF_X1 port map( D => SIG_in_int_23_port, CK => clk, Q 
                           => SIG_in(23), QN => n_1200);
   SIG_in_reg_19_inst : DFF_X1 port map( D => SIG_in_int_19_port, CK => clk, Q 
                           => SIG_in(19), QN => n_1201);
   SIG_in_reg_27_inst : DFF_X1 port map( D => SIG_in_int_27_port, CK => clk, Q 
                           => SIG_in(27), QN => n_1202);
   U3 : AND2_X1 port map( A1 => A_EXP(7), A2 => B_EXP(7), ZN => EXP_pos_int);
   U4 : NAND4_X1 port map( A1 => B_EXP(5), A2 => B_EXP(6), A3 => B_EXP(3), A4 
                           => B_EXP(4), ZN => n4);
   U5 : INV_X1 port map( A => B_EXP(0), ZN => n3);
   U6 : INV_X1 port map( A => B_EXP(2), ZN => n2);
   U7 : INV_X1 port map( A => B_EXP(1), ZN => n1);
   U8 : NOR4_X1 port map( A1 => n4, A2 => n3, A3 => n2, A4 => n1, ZN => n10);
   U9 : NAND4_X1 port map( A1 => A_EXP(5), A2 => A_EXP(6), A3 => A_EXP(3), A4 
                           => A_EXP(4), ZN => n8);
   U10 : INV_X1 port map( A => A_EXP(0), ZN => n7);
   U11 : INV_X1 port map( A => A_EXP(2), ZN => n6);
   U12 : INV_X1 port map( A => A_EXP(1), ZN => n5);
   U13 : NOR4_X1 port map( A1 => n8, A2 => n7, A3 => n6, A4 => n5, ZN => n9);
   U14 : NOR4_X1 port map( A1 => B_EXP(7), A2 => A_EXP(7), A3 => n10, A4 => n9,
                           ZN => N0);
   U15 : INV_X1 port map( A => mw_I4sum_7_port, ZN => n11);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage1 is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         A_EXP : out std_logic_vector (7 downto 0);  A_SIG : out 
         std_logic_vector (31 downto 0);  B_EXP : out std_logic_vector (7 
         downto 0);  B_SIG : out std_logic_vector (31 downto 0);  
         SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : out 
         std_logic);

end FPmul_stage1;

architecture SYN_struct of FPmul_stage1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component UnpackFP_1
      port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector
            (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, 
            isNaN, isINF, isZ, isDN : out std_logic);
   end component;
   
   component UnpackFP_0
      port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector
            (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, 
            isNaN, isINF, isZ, isDN : out std_logic);
   end component;
   
   signal SIGN_out_int, A_EXP_int_7_port, A_EXP_int_6_port, A_EXP_int_5_port, 
      A_EXP_int_4_port, A_EXP_int_3_port, A_EXP_int_2_port, A_EXP_int_1_port, 
      A_EXP_int_0_port, A_SIG_int_23_port, A_SIG_int_22_port, A_SIG_int_21_port
      , A_SIG_int_20_port, A_SIG_int_19_port, A_SIG_int_18_port, 
      A_SIG_int_17_port, A_SIG_int_16_port, A_SIG_int_15_port, 
      A_SIG_int_14_port, A_SIG_int_13_port, A_SIG_int_12_port, 
      A_SIG_int_11_port, A_SIG_int_10_port, A_SIG_int_9_port, A_SIG_int_8_port,
      A_SIG_int_7_port, A_SIG_int_6_port, A_SIG_int_5_port, A_SIG_int_4_port, 
      A_SIG_int_3_port, A_SIG_int_2_port, A_SIG_int_1_port, A_SIG_int_0_port, 
      isINF_int, isNaN_int, isZ_tab_int, B_EXP_int_7_port, B_EXP_int_6_port, 
      B_EXP_int_5_port, B_EXP_int_4_port, B_EXP_int_3_port, B_EXP_int_2_port, 
      B_EXP_int_1_port, B_EXP_int_0_port, B_SIG_int_23_port, B_SIG_int_22_port,
      B_SIG_int_21_port, B_SIG_int_20_port, B_SIG_int_19_port, 
      B_SIG_int_18_port, B_SIG_int_17_port, B_SIG_int_16_port, 
      B_SIG_int_15_port, B_SIG_int_14_port, B_SIG_int_13_port, 
      B_SIG_int_12_port, B_SIG_int_11_port, B_SIG_int_10_port, B_SIG_int_9_port
      , B_SIG_int_8_port, B_SIG_int_7_port, B_SIG_int_6_port, B_SIG_int_5_port,
      B_SIG_int_4_port, B_SIG_int_3_port, B_SIG_int_2_port, B_SIG_int_1_port, 
      B_SIG_int_0_port, A_isINF, A_isNaN, A_isZ, B_isINF, B_isNaN, B_isZ, 
      A_SIGN, B_SIGN, n1, n3, n5, n7, n9, n11, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n_1203, n_1204, n_1205, n_1206, n_1207, 
      n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, 
      n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, 
      n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, 
      n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, 
      n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, 
      n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, 
      n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, 
      n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, 
      n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288 : 
      std_logic;

begin
   
   SIGN_out_stage1_reg : DFF_X1 port map( D => SIGN_out_int, CK => clk, Q => 
                           SIGN_out_stage1, QN => n_1203);
   A_EXP_reg_7_inst : DFF_X1 port map( D => A_EXP_int_7_port, CK => clk, Q => 
                           A_EXP(7), QN => n_1204);
   A_EXP_reg_6_inst : DFF_X1 port map( D => A_EXP_int_6_port, CK => clk, Q => 
                           A_EXP(6), QN => n_1205);
   A_EXP_reg_5_inst : DFF_X1 port map( D => A_EXP_int_5_port, CK => clk, Q => 
                           A_EXP(5), QN => n_1206);
   A_EXP_reg_4_inst : DFF_X1 port map( D => A_EXP_int_4_port, CK => clk, Q => 
                           A_EXP(4), QN => n_1207);
   A_EXP_reg_3_inst : DFF_X1 port map( D => A_EXP_int_3_port, CK => clk, Q => 
                           A_EXP(3), QN => n_1208);
   A_EXP_reg_2_inst : DFF_X1 port map( D => A_EXP_int_2_port, CK => clk, Q => 
                           A_EXP(2), QN => n_1209);
   A_EXP_reg_1_inst : DFF_X1 port map( D => A_EXP_int_1_port, CK => clk, Q => 
                           A_EXP(1), QN => n_1210);
   A_EXP_reg_0_inst : DFF_X1 port map( D => A_EXP_int_0_port, CK => clk, Q => 
                           A_EXP(0), QN => n_1211);
   A_SIG_reg_22_inst : DFF_X1 port map( D => A_SIG_int_22_port, CK => clk, Q =>
                           A_SIG(22), QN => n_1212);
   A_SIG_reg_21_inst : DFF_X1 port map( D => A_SIG_int_21_port, CK => clk, Q =>
                           A_SIG(21), QN => n_1213);
   A_SIG_reg_20_inst : DFF_X1 port map( D => A_SIG_int_20_port, CK => clk, Q =>
                           A_SIG(20), QN => n_1214);
   A_SIG_reg_19_inst : DFF_X1 port map( D => A_SIG_int_19_port, CK => clk, Q =>
                           A_SIG(19), QN => n_1215);
   A_SIG_reg_18_inst : DFF_X1 port map( D => A_SIG_int_18_port, CK => clk, Q =>
                           A_SIG(18), QN => n_1216);
   A_SIG_reg_15_inst : DFF_X1 port map( D => A_SIG_int_15_port, CK => clk, Q =>
                           A_SIG(15), QN => n_1217);
   A_SIG_reg_14_inst : DFF_X1 port map( D => A_SIG_int_14_port, CK => clk, Q =>
                           A_SIG(14), QN => n_1218);
   A_SIG_reg_13_inst : DFF_X1 port map( D => A_SIG_int_13_port, CK => clk, Q =>
                           A_SIG(13), QN => n_1219);
   A_SIG_reg_10_inst : DFF_X1 port map( D => A_SIG_int_10_port, CK => clk, Q =>
                           A_SIG(10), QN => n_1220);
   A_SIG_reg_6_inst : DFF_X1 port map( D => A_SIG_int_6_port, CK => clk, Q => 
                           A_SIG(6), QN => n_1221);
   A_SIG_reg_5_inst : DFF_X1 port map( D => A_SIG_int_5_port, CK => clk, Q => 
                           A_SIG(5), QN => n_1222);
   A_SIG_reg_4_inst : DFF_X1 port map( D => A_SIG_int_4_port, CK => clk, Q => 
                           A_SIG(4), QN => n_1223);
   A_SIG_reg_3_inst : DFF_X1 port map( D => A_SIG_int_3_port, CK => clk, Q => 
                           A_SIG(3), QN => n_1224);
   A_SIG_reg_2_inst : DFF_X1 port map( D => A_SIG_int_2_port, CK => clk, Q => 
                           A_SIG(2), QN => n_1225);
   A_SIG_reg_1_inst : DFF_X1 port map( D => A_SIG_int_1_port, CK => clk, Q => 
                           A_SIG(1), QN => n_1226);
   A_SIG_reg_0_inst : DFF_X1 port map( D => A_SIG_int_0_port, CK => clk, Q => 
                           A_SIG(0), QN => n_1227);
   isINF_stage1_reg : DFF_X1 port map( D => isINF_int, CK => clk, Q => 
                           isINF_stage1, QN => n_1228);
   isNaN_stage1_reg : DFF_X1 port map( D => isNaN_int, CK => clk, Q => 
                           isNaN_stage1, QN => n_1229);
   isZ_tab_stage1_reg : DFF_X1 port map( D => isZ_tab_int, CK => clk, Q => 
                           isZ_tab_stage1, QN => n_1230);
   B_EXP_reg_7_inst : DFF_X1 port map( D => B_EXP_int_7_port, CK => clk, Q => 
                           B_EXP(7), QN => n_1231);
   B_EXP_reg_6_inst : DFF_X1 port map( D => B_EXP_int_6_port, CK => clk, Q => 
                           B_EXP(6), QN => n_1232);
   B_EXP_reg_5_inst : DFF_X1 port map( D => B_EXP_int_5_port, CK => clk, Q => 
                           B_EXP(5), QN => n_1233);
   B_EXP_reg_4_inst : DFF_X1 port map( D => B_EXP_int_4_port, CK => clk, Q => 
                           B_EXP(4), QN => n_1234);
   B_EXP_reg_3_inst : DFF_X1 port map( D => B_EXP_int_3_port, CK => clk, Q => 
                           B_EXP(3), QN => n_1235);
   B_EXP_reg_2_inst : DFF_X1 port map( D => B_EXP_int_2_port, CK => clk, Q => 
                           B_EXP(2), QN => n_1236);
   B_EXP_reg_1_inst : DFF_X1 port map( D => B_EXP_int_1_port, CK => clk, Q => 
                           B_EXP(1), QN => n_1237);
   B_EXP_reg_0_inst : DFF_X1 port map( D => B_EXP_int_0_port, CK => clk, Q => 
                           B_EXP(0), QN => n_1238);
   B_SIG_reg_22_inst : DFF_X1 port map( D => B_SIG_int_22_port, CK => clk, Q =>
                           B_SIG(22), QN => n_1239);
   B_SIG_reg_20_inst : DFF_X1 port map( D => B_SIG_int_20_port, CK => clk, Q =>
                           B_SIG(20), QN => n_1240);
   B_SIG_reg_18_inst : DFF_X1 port map( D => B_SIG_int_18_port, CK => clk, Q =>
                           B_SIG(18), QN => n_1241);
   B_SIG_reg_16_inst : DFF_X1 port map( D => B_SIG_int_16_port, CK => clk, Q =>
                           B_SIG(16), QN => n_1242);
   B_SIG_reg_14_inst : DFF_X1 port map( D => B_SIG_int_14_port, CK => clk, Q =>
                           B_SIG(14), QN => n_1243);
   B_SIG_reg_12_inst : DFF_X1 port map( D => B_SIG_int_12_port, CK => clk, Q =>
                           B_SIG(12), QN => n_1244);
   B_SIG_reg_10_inst : DFF_X1 port map( D => B_SIG_int_10_port, CK => clk, Q =>
                           B_SIG(10), QN => n_1245);
   B_SIG_reg_8_inst : DFF_X1 port map( D => B_SIG_int_8_port, CK => clk, Q => 
                           B_SIG(8), QN => n_1246);
   B_SIG_reg_6_inst : DFF_X1 port map( D => B_SIG_int_6_port, CK => clk, Q => 
                           B_SIG(6), QN => n_1247);
   B_SIG_reg_4_inst : DFF_X1 port map( D => B_SIG_int_4_port, CK => clk, Q => 
                           B_SIG(4), QN => n_1248);
   B_SIG_reg_2_inst : DFF_X1 port map( D => B_SIG_int_2_port, CK => clk, Q => 
                           B_SIG(2), QN => n_1249);
   B_SIG_reg_0_inst : DFF_X1 port map( D => B_SIG_int_0_port, CK => clk, Q => 
                           B_SIG(0), QN => n_1250);
   I0 : UnpackFP_0 port map( FP(31) => FP_A(31), FP(30) => FP_A(30), FP(29) => 
                           FP_A(29), FP(28) => FP_A(28), FP(27) => FP_A(27), 
                           FP(26) => FP_A(26), FP(25) => FP_A(25), FP(24) => 
                           FP_A(24), FP(23) => FP_A(23), FP(22) => FP_A(22), 
                           FP(21) => FP_A(21), FP(20) => FP_A(20), FP(19) => 
                           FP_A(19), FP(18) => FP_A(18), FP(17) => FP_A(17), 
                           FP(16) => FP_A(16), FP(15) => FP_A(15), FP(14) => 
                           FP_A(14), FP(13) => FP_A(13), FP(12) => FP_A(12), 
                           FP(11) => FP_A(11), FP(10) => FP_A(10), FP(9) => 
                           FP_A(9), FP(8) => FP_A(8), FP(7) => FP_A(7), FP(6) 
                           => FP_A(6), FP(5) => FP_A(5), FP(4) => FP_A(4), 
                           FP(3) => FP_A(3), FP(2) => FP_A(2), FP(1) => FP_A(1)
                           , FP(0) => FP_A(0), SIG(31) => n_1251, SIG(30) => 
                           n_1252, SIG(29) => n_1253, SIG(28) => n_1254, 
                           SIG(27) => n_1255, SIG(26) => n_1256, SIG(25) => 
                           n_1257, SIG(24) => n_1258, SIG(23) => 
                           A_SIG_int_23_port, SIG(22) => A_SIG_int_22_port, 
                           SIG(21) => A_SIG_int_21_port, SIG(20) => 
                           A_SIG_int_20_port, SIG(19) => A_SIG_int_19_port, 
                           SIG(18) => A_SIG_int_18_port, SIG(17) => 
                           A_SIG_int_17_port, SIG(16) => A_SIG_int_16_port, 
                           SIG(15) => A_SIG_int_15_port, SIG(14) => 
                           A_SIG_int_14_port, SIG(13) => A_SIG_int_13_port, 
                           SIG(12) => A_SIG_int_12_port, SIG(11) => 
                           A_SIG_int_11_port, SIG(10) => A_SIG_int_10_port, 
                           SIG(9) => A_SIG_int_9_port, SIG(8) => 
                           A_SIG_int_8_port, SIG(7) => A_SIG_int_7_port, SIG(6)
                           => A_SIG_int_6_port, SIG(5) => A_SIG_int_5_port, 
                           SIG(4) => A_SIG_int_4_port, SIG(3) => 
                           A_SIG_int_3_port, SIG(2) => A_SIG_int_2_port, SIG(1)
                           => A_SIG_int_1_port, SIG(0) => A_SIG_int_0_port, 
                           EXP(7) => A_EXP_int_7_port, EXP(6) => 
                           A_EXP_int_6_port, EXP(5) => A_EXP_int_5_port, EXP(4)
                           => A_EXP_int_4_port, EXP(3) => A_EXP_int_3_port, 
                           EXP(2) => A_EXP_int_2_port, EXP(1) => 
                           A_EXP_int_1_port, EXP(0) => A_EXP_int_0_port, SIGN 
                           => A_SIGN, isNaN => A_isNaN, isINF => A_isINF, isZ 
                           => A_isZ, isDN => n_1259);
   I1 : UnpackFP_1 port map( FP(31) => FP_B(31), FP(30) => FP_B(30), FP(29) => 
                           FP_B(29), FP(28) => FP_B(28), FP(27) => FP_B(27), 
                           FP(26) => FP_B(26), FP(25) => FP_B(25), FP(24) => 
                           FP_B(24), FP(23) => FP_B(23), FP(22) => FP_B(22), 
                           FP(21) => FP_B(21), FP(20) => FP_B(20), FP(19) => 
                           FP_B(19), FP(18) => FP_B(18), FP(17) => FP_B(17), 
                           FP(16) => FP_B(16), FP(15) => FP_B(15), FP(14) => 
                           FP_B(14), FP(13) => FP_B(13), FP(12) => FP_B(12), 
                           FP(11) => FP_B(11), FP(10) => FP_B(10), FP(9) => 
                           FP_B(9), FP(8) => FP_B(8), FP(7) => FP_B(7), FP(6) 
                           => FP_B(6), FP(5) => FP_B(5), FP(4) => FP_B(4), 
                           FP(3) => FP_B(3), FP(2) => FP_B(2), FP(1) => FP_B(1)
                           , FP(0) => FP_B(0), SIG(31) => n_1260, SIG(30) => 
                           n_1261, SIG(29) => n_1262, SIG(28) => n_1263, 
                           SIG(27) => n_1264, SIG(26) => n_1265, SIG(25) => 
                           n_1266, SIG(24) => n_1267, SIG(23) => 
                           B_SIG_int_23_port, SIG(22) => B_SIG_int_22_port, 
                           SIG(21) => B_SIG_int_21_port, SIG(20) => 
                           B_SIG_int_20_port, SIG(19) => B_SIG_int_19_port, 
                           SIG(18) => B_SIG_int_18_port, SIG(17) => 
                           B_SIG_int_17_port, SIG(16) => B_SIG_int_16_port, 
                           SIG(15) => B_SIG_int_15_port, SIG(14) => 
                           B_SIG_int_14_port, SIG(13) => B_SIG_int_13_port, 
                           SIG(12) => B_SIG_int_12_port, SIG(11) => 
                           B_SIG_int_11_port, SIG(10) => B_SIG_int_10_port, 
                           SIG(9) => B_SIG_int_9_port, SIG(8) => 
                           B_SIG_int_8_port, SIG(7) => B_SIG_int_7_port, SIG(6)
                           => B_SIG_int_6_port, SIG(5) => B_SIG_int_5_port, 
                           SIG(4) => B_SIG_int_4_port, SIG(3) => 
                           B_SIG_int_3_port, SIG(2) => B_SIG_int_2_port, SIG(1)
                           => B_SIG_int_1_port, SIG(0) => B_SIG_int_0_port, 
                           EXP(7) => B_EXP_int_7_port, EXP(6) => 
                           B_EXP_int_6_port, EXP(5) => B_EXP_int_5_port, EXP(4)
                           => B_EXP_int_4_port, EXP(3) => B_EXP_int_3_port, 
                           EXP(2) => B_EXP_int_2_port, EXP(1) => 
                           B_EXP_int_1_port, EXP(0) => B_EXP_int_0_port, SIGN 
                           => B_SIGN, isNaN => B_isNaN, isINF => B_isINF, isZ 
                           => B_isZ, isDN => n_1268);
   A_SIG_reg_9_inst : DFF_X1 port map( D => A_SIG_int_9_port, CK => clk, Q => 
                           A_SIG(9), QN => n_1269);
   A_SIG_reg_7_inst : DFF_X1 port map( D => A_SIG_int_7_port, CK => clk, Q => 
                           A_SIG(7), QN => n_1270);
   A_SIG_reg_8_inst : DFF_X1 port map( D => A_SIG_int_8_port, CK => clk, Q => 
                           A_SIG(8), QN => n_1271);
   A_SIG_reg_11_inst : DFF_X1 port map( D => A_SIG_int_11_port, CK => clk, Q =>
                           A_SIG(11), QN => n_1272);
   A_SIG_reg_17_inst : DFF_X1 port map( D => A_SIG_int_17_port, CK => clk, Q =>
                           A_SIG(17), QN => n_1273);
   A_SIG_reg_16_inst : DFF_X1 port map( D => A_SIG_int_16_port, CK => clk, Q =>
                           A_SIG(16), QN => n_1274);
   A_SIG_reg_12_inst : DFF_X1 port map( D => A_SIG_int_12_port, CK => clk, Q =>
                           A_SIG(12), QN => n_1275);
   A_SIG_reg_23_inst : DFF_X1 port map( D => A_SIG_int_23_port, CK => clk, Q =>
                           A_SIG(23), QN => n_1276);
   B_SIG_reg_23_inst : DFF_X1 port map( D => B_SIG_int_23_port, CK => clk, Q =>
                           B_SIG(23), QN => n_1277);
   B_SIG_reg_1_inst : SDFF_X1 port map( D => B_SIG_int_1_port, SI => n11, SE =>
                           n11, CK => clk, Q => B_SIG(1), QN => n_1278);
   B_SIG_reg_19_inst : DFF_X2 port map( D => B_SIG_int_19_port, CK => clk, Q =>
                           B_SIG(19), QN => n_1279);
   B_SIG_reg_11_inst : DFF_X2 port map( D => B_SIG_int_11_port, CK => clk, Q =>
                           B_SIG(11), QN => n_1280);
   B_SIG_reg_5_inst : DFF_X2 port map( D => B_SIG_int_5_port, CK => clk, Q => 
                           B_SIG(5), QN => n_1281);
   B_SIG_reg_3_inst : DFF_X1 port map( D => B_SIG_int_3_port, CK => clk, Q => 
                           n_1282, QN => n9);
   B_SIG_reg_21_inst : DFF_X1 port map( D => B_SIG_int_21_port, CK => clk, Q =>
                           n_1283, QN => n7);
   B_SIG_reg_7_inst : DFF_X1 port map( D => B_SIG_int_7_port, CK => clk, Q => 
                           n_1284, QN => n5);
   B_SIG_reg_9_inst : DFF_X2 port map( D => B_SIG_int_9_port, CK => clk, Q => 
                           B_SIG(9), QN => n_1285);
   B_SIG_reg_15_inst : DFF_X1 port map( D => B_SIG_int_15_port, CK => clk, Q =>
                           n_1286, QN => n3);
   B_SIG_reg_13_inst : DFF_X1 port map( D => B_SIG_int_13_port, CK => clk, Q =>
                           n_1287, QN => n1);
   B_SIG_reg_17_inst : DFF_X2 port map( D => B_SIG_int_17_port, CK => clk, Q =>
                           B_SIG(17), QN => n_1288);
   U3 : INV_X2 port map( A => n1, ZN => B_SIG(13));
   U4 : INV_X2 port map( A => n3, ZN => B_SIG(15));
   U5 : INV_X2 port map( A => n5, ZN => B_SIG(7));
   U6 : INV_X2 port map( A => n7, ZN => B_SIG(21));
   U7 : INV_X2 port map( A => n9, ZN => B_SIG(3));
   n11 <= '0';
   A_SIG(31) <= '0';
   A_SIG(30) <= '0';
   A_SIG(29) <= '0';
   A_SIG(28) <= '0';
   A_SIG(27) <= '0';
   A_SIG(26) <= '0';
   A_SIG(25) <= '0';
   A_SIG(24) <= '0';
   B_SIG(31) <= '0';
   B_SIG(30) <= '0';
   B_SIG(28) <= '0';
   B_SIG(27) <= '0';
   B_SIG(26) <= '0';
   B_SIG(25) <= '0';
   B_SIG(24) <= '0';
   B_SIG(29) <= '0';
   U25 : INV_X1 port map( A => B_isZ, ZN => n20);
   U26 : INV_X1 port map( A => A_isZ, ZN => n22);
   U27 : OR2_X1 port map( A1 => B_isNaN, A2 => A_isNaN, ZN => n21);
   U28 : INV_X1 port map( A => n21, ZN => n18);
   U29 : INV_X1 port map( A => A_isINF, ZN => n25);
   U30 : NAND2_X1 port map( A1 => n18, A2 => n25, ZN => n19);
   U31 : AOI211_X1 port map( C1 => n20, C2 => n22, A => n19, B => B_isINF, ZN 
                           => isZ_tab_int);
   U32 : NAND2_X1 port map( A1 => B_isZ, A2 => A_isINF, ZN => n26);
   U33 : NAND2_X1 port map( A1 => n21, A2 => n25, ZN => n23);
   U34 : MUX2_X1 port map( A => n23, B => n22, S => B_isINF, Z => n24);
   U35 : NAND2_X1 port map( A1 => n26, A2 => n24, ZN => isNaN_int);
   U36 : NOR2_X1 port map( A1 => B_isZ, A2 => n25, ZN => n29);
   U37 : INV_X1 port map( A => n26, ZN => n27);
   U38 : NOR2_X1 port map( A1 => A_isZ, A2 => n27, ZN => n28);
   U39 : MUX2_X1 port map( A => n29, B => n28, S => B_isINF, Z => isINF_int);
   U40 : XOR2_X1 port map( A => B_SIGN, B => A_SIGN, Z => SIGN_out_int);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         FP_Z : out std_logic_vector (31 downto 0));

end FPmul;

architecture SYN_pipeline of FPmul is

   component FPmul_stage4
      port( EXP_neg : in std_logic;  EXP_out_round : in std_logic_vector (7 
            downto 0);  EXP_pos, SIGN_out : in std_logic;  SIG_out_round : in 
            std_logic_vector (27 downto 0);  clk, isINF_tab, isNaN, isZ_tab : 
            in std_logic;  FP_Z : out std_logic_vector (31 downto 0));
   end component;
   
   component FPmul_stage3
      port( EXP_in : in std_logic_vector (7 downto 0);  EXP_neg_stage2, 
            EXP_pos_stage2, SIGN_out_stage2 : in std_logic;  SIG_in : in 
            std_logic_vector (27 downto 0);  clk, isINF_stage2, isNaN_stage2, 
            isZ_tab_stage2 : in std_logic;  EXP_neg : out std_logic;  
            EXP_out_round : out std_logic_vector (7 downto 0);  EXP_pos, 
            SIGN_out : out std_logic;  SIG_out_round : out std_logic_vector (27
            downto 0);  isINF_tab, isNaN, isZ_tab : out std_logic);
   end component;
   
   component FPmul_stage2
      port( A_EXP : in std_logic_vector (7 downto 0);  A_SIG : in 
            std_logic_vector (31 downto 0);  B_EXP : in std_logic_vector (7 
            downto 0);  B_SIG : in std_logic_vector (31 downto 0);  
            SIGN_out_stage1, clk, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : 
            in std_logic;  EXP_in : out std_logic_vector (7 downto 0);  
            EXP_neg_stage2, EXP_pos_stage2, SIGN_out_stage2 : out std_logic;  
            SIG_in : out std_logic_vector (27 downto 0);  isINF_stage2, 
            isNaN_stage2, isZ_tab_stage2 : out std_logic);
   end component;
   
   component FPmul_stage1
      port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic
            ;  A_EXP : out std_logic_vector (7 downto 0);  A_SIG : out 
            std_logic_vector (31 downto 0);  B_EXP : out std_logic_vector (7 
            downto 0);  B_SIG : out std_logic_vector (31 downto 0);  
            SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : out 
            std_logic);
   end component;
   
   signal A_EXP_7_port, A_EXP_6_port, A_EXP_5_port, A_EXP_4_port, A_EXP_3_port,
      A_EXP_2_port, A_EXP_1_port, A_EXP_0_port, A_SIG_23_port, A_SIG_22_port, 
      A_SIG_21_port, A_SIG_20_port, A_SIG_19_port, A_SIG_18_port, A_SIG_17_port
      , A_SIG_16_port, A_SIG_15_port, A_SIG_14_port, A_SIG_13_port, 
      A_SIG_12_port, A_SIG_11_port, A_SIG_10_port, A_SIG_9_port, A_SIG_8_port, 
      A_SIG_7_port, A_SIG_6_port, A_SIG_5_port, A_SIG_4_port, A_SIG_3_port, 
      A_SIG_2_port, A_SIG_1_port, A_SIG_0_port, B_EXP_7_port, B_EXP_6_port, 
      B_EXP_5_port, B_EXP_4_port, B_EXP_3_port, B_EXP_2_port, B_EXP_1_port, 
      B_EXP_0_port, B_SIG_23_port, B_SIG_22_port, B_SIG_21_port, B_SIG_20_port,
      B_SIG_19_port, B_SIG_18_port, B_SIG_17_port, B_SIG_16_port, B_SIG_15_port
      , B_SIG_14_port, B_SIG_13_port, B_SIG_12_port, B_SIG_11_port, 
      B_SIG_10_port, B_SIG_9_port, B_SIG_8_port, B_SIG_7_port, B_SIG_6_port, 
      B_SIG_5_port, B_SIG_4_port, B_SIG_3_port, B_SIG_2_port, B_SIG_1_port, 
      B_SIG_0_port, SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1
      , EXP_in_7_port, EXP_in_6_port, EXP_in_5_port, EXP_in_4_port, 
      EXP_in_3_port, EXP_in_2_port, EXP_in_1_port, EXP_in_0_port, 
      EXP_neg_stage2, EXP_pos_stage2, SIGN_out_stage2, SIG_in_27_port, 
      SIG_in_26_port, SIG_in_25_port, SIG_in_24_port, SIG_in_23_port, 
      SIG_in_22_port, SIG_in_21_port, SIG_in_20_port, SIG_in_19_port, 
      SIG_in_18_port, SIG_in_17_port, SIG_in_16_port, SIG_in_15_port, 
      SIG_in_14_port, SIG_in_13_port, SIG_in_12_port, SIG_in_11_port, 
      SIG_in_10_port, SIG_in_9_port, SIG_in_8_port, SIG_in_7_port, 
      SIG_in_6_port, SIG_in_5_port, SIG_in_4_port, SIG_in_3_port, SIG_in_2_port
      , SIG_in_1_port, SIG_in_0_port, isINF_stage2, isNaN_stage2, 
      isZ_tab_stage2, EXP_neg, EXP_out_round_7_port, EXP_out_round_6_port, 
      EXP_out_round_5_port, EXP_out_round_4_port, EXP_out_round_3_port, 
      EXP_out_round_2_port, EXP_out_round_1_port, EXP_out_round_0_port, EXP_pos
      , SIGN_out, SIG_out_round_27_port, SIG_out_round_26_port, 
      SIG_out_round_25_port, SIG_out_round_24_port, SIG_out_round_23_port, 
      SIG_out_round_22_port, SIG_out_round_21_port, SIG_out_round_20_port, 
      SIG_out_round_19_port, SIG_out_round_18_port, SIG_out_round_17_port, 
      SIG_out_round_16_port, SIG_out_round_15_port, SIG_out_round_14_port, 
      SIG_out_round_13_port, SIG_out_round_12_port, SIG_out_round_11_port, 
      SIG_out_round_10_port, SIG_out_round_9_port, SIG_out_round_8_port, 
      SIG_out_round_7_port, SIG_out_round_6_port, SIG_out_round_5_port, 
      SIG_out_round_4_port, SIG_out_round_3_port, SIG_out_round_1_port, 
      SIG_out_round_0_port, isINF_tab, isNaN, isZ_tab, n1, n_1289, n_1290, 
      n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, 
      n_1300, n_1301, n_1302, n_1303, n_1304, n_1305 : std_logic;

begin
   
   I1 : FPmul_stage1 port map( FP_A(31) => FP_A(31), FP_A(30) => FP_A(30), 
                           FP_A(29) => FP_A(29), FP_A(28) => FP_A(28), FP_A(27)
                           => FP_A(27), FP_A(26) => FP_A(26), FP_A(25) => 
                           FP_A(25), FP_A(24) => FP_A(24), FP_A(23) => FP_A(23)
                           , FP_A(22) => FP_A(22), FP_A(21) => FP_A(21), 
                           FP_A(20) => FP_A(20), FP_A(19) => FP_A(19), FP_A(18)
                           => FP_A(18), FP_A(17) => FP_A(17), FP_A(16) => 
                           FP_A(16), FP_A(15) => FP_A(15), FP_A(14) => FP_A(14)
                           , FP_A(13) => FP_A(13), FP_A(12) => FP_A(12), 
                           FP_A(11) => FP_A(11), FP_A(10) => FP_A(10), FP_A(9) 
                           => FP_A(9), FP_A(8) => FP_A(8), FP_A(7) => FP_A(7), 
                           FP_A(6) => FP_A(6), FP_A(5) => FP_A(5), FP_A(4) => 
                           FP_A(4), FP_A(3) => FP_A(3), FP_A(2) => FP_A(2), 
                           FP_A(1) => FP_A(1), FP_A(0) => FP_A(0), FP_B(31) => 
                           FP_B(31), FP_B(30) => FP_B(30), FP_B(29) => FP_B(29)
                           , FP_B(28) => FP_B(28), FP_B(27) => FP_B(27), 
                           FP_B(26) => FP_B(26), FP_B(25) => FP_B(25), FP_B(24)
                           => FP_B(24), FP_B(23) => FP_B(23), FP_B(22) => 
                           FP_B(22), FP_B(21) => FP_B(21), FP_B(20) => FP_B(20)
                           , FP_B(19) => FP_B(19), FP_B(18) => FP_B(18), 
                           FP_B(17) => FP_B(17), FP_B(16) => FP_B(16), FP_B(15)
                           => FP_B(15), FP_B(14) => FP_B(14), FP_B(13) => 
                           FP_B(13), FP_B(12) => FP_B(12), FP_B(11) => FP_B(11)
                           , FP_B(10) => FP_B(10), FP_B(9) => FP_B(9), FP_B(8) 
                           => FP_B(8), FP_B(7) => FP_B(7), FP_B(6) => FP_B(6), 
                           FP_B(5) => FP_B(5), FP_B(4) => FP_B(4), FP_B(3) => 
                           FP_B(3), FP_B(2) => FP_B(2), FP_B(1) => FP_B(1), 
                           FP_B(0) => FP_B(0), clk => clk, A_EXP(7) => 
                           A_EXP_7_port, A_EXP(6) => A_EXP_6_port, A_EXP(5) => 
                           A_EXP_5_port, A_EXP(4) => A_EXP_4_port, A_EXP(3) => 
                           A_EXP_3_port, A_EXP(2) => A_EXP_2_port, A_EXP(1) => 
                           A_EXP_1_port, A_EXP(0) => A_EXP_0_port, A_SIG(31) =>
                           n_1289, A_SIG(30) => n_1290, A_SIG(29) => n_1291, 
                           A_SIG(28) => n_1292, A_SIG(27) => n_1293, A_SIG(26) 
                           => n_1294, A_SIG(25) => n_1295, A_SIG(24) => n_1296,
                           A_SIG(23) => A_SIG_23_port, A_SIG(22) => 
                           A_SIG_22_port, A_SIG(21) => A_SIG_21_port, A_SIG(20)
                           => A_SIG_20_port, A_SIG(19) => A_SIG_19_port, 
                           A_SIG(18) => A_SIG_18_port, A_SIG(17) => 
                           A_SIG_17_port, A_SIG(16) => A_SIG_16_port, A_SIG(15)
                           => A_SIG_15_port, A_SIG(14) => A_SIG_14_port, 
                           A_SIG(13) => A_SIG_13_port, A_SIG(12) => 
                           A_SIG_12_port, A_SIG(11) => A_SIG_11_port, A_SIG(10)
                           => A_SIG_10_port, A_SIG(9) => A_SIG_9_port, A_SIG(8)
                           => A_SIG_8_port, A_SIG(7) => A_SIG_7_port, A_SIG(6) 
                           => A_SIG_6_port, A_SIG(5) => A_SIG_5_port, A_SIG(4) 
                           => A_SIG_4_port, A_SIG(3) => A_SIG_3_port, A_SIG(2) 
                           => A_SIG_2_port, A_SIG(1) => A_SIG_1_port, A_SIG(0) 
                           => A_SIG_0_port, B_EXP(7) => B_EXP_7_port, B_EXP(6) 
                           => B_EXP_6_port, B_EXP(5) => B_EXP_5_port, B_EXP(4) 
                           => B_EXP_4_port, B_EXP(3) => B_EXP_3_port, B_EXP(2) 
                           => B_EXP_2_port, B_EXP(1) => B_EXP_1_port, B_EXP(0) 
                           => B_EXP_0_port, B_SIG(31) => n_1297, B_SIG(30) => 
                           n_1298, B_SIG(29) => n_1299, B_SIG(28) => n_1300, 
                           B_SIG(27) => n_1301, B_SIG(26) => n_1302, B_SIG(25) 
                           => n_1303, B_SIG(24) => n_1304, B_SIG(23) => 
                           B_SIG_23_port, B_SIG(22) => B_SIG_22_port, B_SIG(21)
                           => B_SIG_21_port, B_SIG(20) => B_SIG_20_port, 
                           B_SIG(19) => B_SIG_19_port, B_SIG(18) => 
                           B_SIG_18_port, B_SIG(17) => B_SIG_17_port, B_SIG(16)
                           => B_SIG_16_port, B_SIG(15) => B_SIG_15_port, 
                           B_SIG(14) => B_SIG_14_port, B_SIG(13) => 
                           B_SIG_13_port, B_SIG(12) => B_SIG_12_port, B_SIG(11)
                           => B_SIG_11_port, B_SIG(10) => B_SIG_10_port, 
                           B_SIG(9) => B_SIG_9_port, B_SIG(8) => B_SIG_8_port, 
                           B_SIG(7) => B_SIG_7_port, B_SIG(6) => B_SIG_6_port, 
                           B_SIG(5) => B_SIG_5_port, B_SIG(4) => B_SIG_4_port, 
                           B_SIG(3) => B_SIG_3_port, B_SIG(2) => B_SIG_2_port, 
                           B_SIG(1) => B_SIG_1_port, B_SIG(0) => B_SIG_0_port, 
                           SIGN_out_stage1 => SIGN_out_stage1, isINF_stage1 => 
                           isINF_stage1, isNaN_stage1 => isNaN_stage1, 
                           isZ_tab_stage1 => isZ_tab_stage1);
   I2 : FPmul_stage2 port map( A_EXP(7) => A_EXP_7_port, A_EXP(6) => 
                           A_EXP_6_port, A_EXP(5) => A_EXP_5_port, A_EXP(4) => 
                           A_EXP_4_port, A_EXP(3) => A_EXP_3_port, A_EXP(2) => 
                           A_EXP_2_port, A_EXP(1) => A_EXP_1_port, A_EXP(0) => 
                           A_EXP_0_port, A_SIG(31) => n1, A_SIG(30) => n1, 
                           A_SIG(29) => n1, A_SIG(28) => n1, A_SIG(27) => n1, 
                           A_SIG(26) => n1, A_SIG(25) => n1, A_SIG(24) => n1, 
                           A_SIG(23) => A_SIG_23_port, A_SIG(22) => 
                           A_SIG_22_port, A_SIG(21) => A_SIG_21_port, A_SIG(20)
                           => A_SIG_20_port, A_SIG(19) => A_SIG_19_port, 
                           A_SIG(18) => A_SIG_18_port, A_SIG(17) => 
                           A_SIG_17_port, A_SIG(16) => A_SIG_16_port, A_SIG(15)
                           => A_SIG_15_port, A_SIG(14) => A_SIG_14_port, 
                           A_SIG(13) => A_SIG_13_port, A_SIG(12) => 
                           A_SIG_12_port, A_SIG(11) => A_SIG_11_port, A_SIG(10)
                           => A_SIG_10_port, A_SIG(9) => A_SIG_9_port, A_SIG(8)
                           => A_SIG_8_port, A_SIG(7) => A_SIG_7_port, A_SIG(6) 
                           => A_SIG_6_port, A_SIG(5) => A_SIG_5_port, A_SIG(4) 
                           => A_SIG_4_port, A_SIG(3) => A_SIG_3_port, A_SIG(2) 
                           => A_SIG_2_port, A_SIG(1) => A_SIG_1_port, A_SIG(0) 
                           => A_SIG_0_port, B_EXP(7) => B_EXP_7_port, B_EXP(6) 
                           => B_EXP_6_port, B_EXP(5) => B_EXP_5_port, B_EXP(4) 
                           => B_EXP_4_port, B_EXP(3) => B_EXP_3_port, B_EXP(2) 
                           => B_EXP_2_port, B_EXP(1) => B_EXP_1_port, B_EXP(0) 
                           => B_EXP_0_port, B_SIG(31) => n1, B_SIG(30) => n1, 
                           B_SIG(29) => n1, B_SIG(28) => n1, B_SIG(27) => n1, 
                           B_SIG(26) => n1, B_SIG(25) => n1, B_SIG(24) => n1, 
                           B_SIG(23) => B_SIG_23_port, B_SIG(22) => 
                           B_SIG_22_port, B_SIG(21) => B_SIG_21_port, B_SIG(20)
                           => B_SIG_20_port, B_SIG(19) => B_SIG_19_port, 
                           B_SIG(18) => B_SIG_18_port, B_SIG(17) => 
                           B_SIG_17_port, B_SIG(16) => B_SIG_16_port, B_SIG(15)
                           => B_SIG_15_port, B_SIG(14) => B_SIG_14_port, 
                           B_SIG(13) => B_SIG_13_port, B_SIG(12) => 
                           B_SIG_12_port, B_SIG(11) => B_SIG_11_port, B_SIG(10)
                           => B_SIG_10_port, B_SIG(9) => B_SIG_9_port, B_SIG(8)
                           => B_SIG_8_port, B_SIG(7) => B_SIG_7_port, B_SIG(6) 
                           => B_SIG_6_port, B_SIG(5) => B_SIG_5_port, B_SIG(4) 
                           => B_SIG_4_port, B_SIG(3) => B_SIG_3_port, B_SIG(2) 
                           => B_SIG_2_port, B_SIG(1) => B_SIG_1_port, B_SIG(0) 
                           => B_SIG_0_port, SIGN_out_stage1 => SIGN_out_stage1,
                           clk => clk, isINF_stage1 => isINF_stage1, 
                           isNaN_stage1 => isNaN_stage1, isZ_tab_stage1 => 
                           isZ_tab_stage1, EXP_in(7) => EXP_in_7_port, 
                           EXP_in(6) => EXP_in_6_port, EXP_in(5) => 
                           EXP_in_5_port, EXP_in(4) => EXP_in_4_port, EXP_in(3)
                           => EXP_in_3_port, EXP_in(2) => EXP_in_2_port, 
                           EXP_in(1) => EXP_in_1_port, EXP_in(0) => 
                           EXP_in_0_port, EXP_neg_stage2 => EXP_neg_stage2, 
                           EXP_pos_stage2 => EXP_pos_stage2, SIGN_out_stage2 =>
                           SIGN_out_stage2, SIG_in(27) => SIG_in_27_port, 
                           SIG_in(26) => SIG_in_26_port, SIG_in(25) => 
                           SIG_in_25_port, SIG_in(24) => SIG_in_24_port, 
                           SIG_in(23) => SIG_in_23_port, SIG_in(22) => 
                           SIG_in_22_port, SIG_in(21) => SIG_in_21_port, 
                           SIG_in(20) => SIG_in_20_port, SIG_in(19) => 
                           SIG_in_19_port, SIG_in(18) => SIG_in_18_port, 
                           SIG_in(17) => SIG_in_17_port, SIG_in(16) => 
                           SIG_in_16_port, SIG_in(15) => SIG_in_15_port, 
                           SIG_in(14) => SIG_in_14_port, SIG_in(13) => 
                           SIG_in_13_port, SIG_in(12) => SIG_in_12_port, 
                           SIG_in(11) => SIG_in_11_port, SIG_in(10) => 
                           SIG_in_10_port, SIG_in(9) => SIG_in_9_port, 
                           SIG_in(8) => SIG_in_8_port, SIG_in(7) => 
                           SIG_in_7_port, SIG_in(6) => SIG_in_6_port, SIG_in(5)
                           => SIG_in_5_port, SIG_in(4) => SIG_in_4_port, 
                           SIG_in(3) => SIG_in_3_port, SIG_in(2) => 
                           SIG_in_2_port, SIG_in(1) => SIG_in_1_port, SIG_in(0)
                           => SIG_in_0_port, isINF_stage2 => isINF_stage2, 
                           isNaN_stage2 => isNaN_stage2, isZ_tab_stage2 => 
                           isZ_tab_stage2);
   I3 : FPmul_stage3 port map( EXP_in(7) => EXP_in_7_port, EXP_in(6) => 
                           EXP_in_6_port, EXP_in(5) => EXP_in_5_port, EXP_in(4)
                           => EXP_in_4_port, EXP_in(3) => EXP_in_3_port, 
                           EXP_in(2) => EXP_in_2_port, EXP_in(1) => 
                           EXP_in_1_port, EXP_in(0) => EXP_in_0_port, 
                           EXP_neg_stage2 => EXP_neg_stage2, EXP_pos_stage2 => 
                           EXP_pos_stage2, SIGN_out_stage2 => SIGN_out_stage2, 
                           SIG_in(27) => SIG_in_27_port, SIG_in(26) => 
                           SIG_in_26_port, SIG_in(25) => SIG_in_25_port, 
                           SIG_in(24) => SIG_in_24_port, SIG_in(23) => 
                           SIG_in_23_port, SIG_in(22) => SIG_in_22_port, 
                           SIG_in(21) => SIG_in_21_port, SIG_in(20) => 
                           SIG_in_20_port, SIG_in(19) => SIG_in_19_port, 
                           SIG_in(18) => SIG_in_18_port, SIG_in(17) => 
                           SIG_in_17_port, SIG_in(16) => SIG_in_16_port, 
                           SIG_in(15) => SIG_in_15_port, SIG_in(14) => 
                           SIG_in_14_port, SIG_in(13) => SIG_in_13_port, 
                           SIG_in(12) => SIG_in_12_port, SIG_in(11) => 
                           SIG_in_11_port, SIG_in(10) => SIG_in_10_port, 
                           SIG_in(9) => SIG_in_9_port, SIG_in(8) => 
                           SIG_in_8_port, SIG_in(7) => SIG_in_7_port, SIG_in(6)
                           => SIG_in_6_port, SIG_in(5) => SIG_in_5_port, 
                           SIG_in(4) => SIG_in_4_port, SIG_in(3) => 
                           SIG_in_3_port, SIG_in(2) => SIG_in_2_port, SIG_in(1)
                           => SIG_in_1_port, SIG_in(0) => SIG_in_0_port, clk =>
                           clk, isINF_stage2 => isINF_stage2, isNaN_stage2 => 
                           isNaN_stage2, isZ_tab_stage2 => isZ_tab_stage2, 
                           EXP_neg => EXP_neg, EXP_out_round(7) => 
                           EXP_out_round_7_port, EXP_out_round(6) => 
                           EXP_out_round_6_port, EXP_out_round(5) => 
                           EXP_out_round_5_port, EXP_out_round(4) => 
                           EXP_out_round_4_port, EXP_out_round(3) => 
                           EXP_out_round_3_port, EXP_out_round(2) => 
                           EXP_out_round_2_port, EXP_out_round(1) => 
                           EXP_out_round_1_port, EXP_out_round(0) => 
                           EXP_out_round_0_port, EXP_pos => EXP_pos, SIGN_out 
                           => SIGN_out, SIG_out_round(27) => 
                           SIG_out_round_27_port, SIG_out_round(26) => 
                           SIG_out_round_26_port, SIG_out_round(25) => 
                           SIG_out_round_25_port, SIG_out_round(24) => 
                           SIG_out_round_24_port, SIG_out_round(23) => 
                           SIG_out_round_23_port, SIG_out_round(22) => 
                           SIG_out_round_22_port, SIG_out_round(21) => 
                           SIG_out_round_21_port, SIG_out_round(20) => 
                           SIG_out_round_20_port, SIG_out_round(19) => 
                           SIG_out_round_19_port, SIG_out_round(18) => 
                           SIG_out_round_18_port, SIG_out_round(17) => 
                           SIG_out_round_17_port, SIG_out_round(16) => 
                           SIG_out_round_16_port, SIG_out_round(15) => 
                           SIG_out_round_15_port, SIG_out_round(14) => 
                           SIG_out_round_14_port, SIG_out_round(13) => 
                           SIG_out_round_13_port, SIG_out_round(12) => 
                           SIG_out_round_12_port, SIG_out_round(11) => 
                           SIG_out_round_11_port, SIG_out_round(10) => 
                           SIG_out_round_10_port, SIG_out_round(9) => 
                           SIG_out_round_9_port, SIG_out_round(8) => 
                           SIG_out_round_8_port, SIG_out_round(7) => 
                           SIG_out_round_7_port, SIG_out_round(6) => 
                           SIG_out_round_6_port, SIG_out_round(5) => 
                           SIG_out_round_5_port, SIG_out_round(4) => 
                           SIG_out_round_4_port, SIG_out_round(3) => 
                           SIG_out_round_3_port, SIG_out_round(2) => n_1305, 
                           SIG_out_round(1) => SIG_out_round_1_port, 
                           SIG_out_round(0) => SIG_out_round_0_port, isINF_tab 
                           => isINF_tab, isNaN => isNaN, isZ_tab => isZ_tab);
   I4 : FPmul_stage4 port map( EXP_neg => EXP_neg, EXP_out_round(7) => 
                           EXP_out_round_7_port, EXP_out_round(6) => 
                           EXP_out_round_6_port, EXP_out_round(5) => 
                           EXP_out_round_5_port, EXP_out_round(4) => 
                           EXP_out_round_4_port, EXP_out_round(3) => 
                           EXP_out_round_3_port, EXP_out_round(2) => 
                           EXP_out_round_2_port, EXP_out_round(1) => 
                           EXP_out_round_1_port, EXP_out_round(0) => 
                           EXP_out_round_0_port, EXP_pos => EXP_pos, SIGN_out 
                           => SIGN_out, SIG_out_round(27) => 
                           SIG_out_round_27_port, SIG_out_round(26) => 
                           SIG_out_round_26_port, SIG_out_round(25) => 
                           SIG_out_round_25_port, SIG_out_round(24) => 
                           SIG_out_round_24_port, SIG_out_round(23) => 
                           SIG_out_round_23_port, SIG_out_round(22) => 
                           SIG_out_round_22_port, SIG_out_round(21) => 
                           SIG_out_round_21_port, SIG_out_round(20) => 
                           SIG_out_round_20_port, SIG_out_round(19) => 
                           SIG_out_round_19_port, SIG_out_round(18) => 
                           SIG_out_round_18_port, SIG_out_round(17) => 
                           SIG_out_round_17_port, SIG_out_round(16) => 
                           SIG_out_round_16_port, SIG_out_round(15) => 
                           SIG_out_round_15_port, SIG_out_round(14) => 
                           SIG_out_round_14_port, SIG_out_round(13) => 
                           SIG_out_round_13_port, SIG_out_round(12) => 
                           SIG_out_round_12_port, SIG_out_round(11) => 
                           SIG_out_round_11_port, SIG_out_round(10) => 
                           SIG_out_round_10_port, SIG_out_round(9) => 
                           SIG_out_round_9_port, SIG_out_round(8) => 
                           SIG_out_round_8_port, SIG_out_round(7) => 
                           SIG_out_round_7_port, SIG_out_round(6) => 
                           SIG_out_round_6_port, SIG_out_round(5) => 
                           SIG_out_round_5_port, SIG_out_round(4) => 
                           SIG_out_round_4_port, SIG_out_round(3) => 
                           SIG_out_round_3_port, SIG_out_round(2) => n1, 
                           SIG_out_round(1) => SIG_out_round_1_port, 
                           SIG_out_round(0) => SIG_out_round_0_port, clk => clk
                           , isINF_tab => isINF_tab, isNaN => isNaN, isZ_tab =>
                           isZ_tab, FP_Z(31) => FP_Z(31), FP_Z(30) => FP_Z(30),
                           FP_Z(29) => FP_Z(29), FP_Z(28) => FP_Z(28), FP_Z(27)
                           => FP_Z(27), FP_Z(26) => FP_Z(26), FP_Z(25) => 
                           FP_Z(25), FP_Z(24) => FP_Z(24), FP_Z(23) => FP_Z(23)
                           , FP_Z(22) => FP_Z(22), FP_Z(21) => FP_Z(21), 
                           FP_Z(20) => FP_Z(20), FP_Z(19) => FP_Z(19), FP_Z(18)
                           => FP_Z(18), FP_Z(17) => FP_Z(17), FP_Z(16) => 
                           FP_Z(16), FP_Z(15) => FP_Z(15), FP_Z(14) => FP_Z(14)
                           , FP_Z(13) => FP_Z(13), FP_Z(12) => FP_Z(12), 
                           FP_Z(11) => FP_Z(11), FP_Z(10) => FP_Z(10), FP_Z(9) 
                           => FP_Z(9), FP_Z(8) => FP_Z(8), FP_Z(7) => FP_Z(7), 
                           FP_Z(6) => FP_Z(6), FP_Z(5) => FP_Z(5), FP_Z(4) => 
                           FP_Z(4), FP_Z(3) => FP_Z(3), FP_Z(2) => FP_Z(2), 
                           FP_Z(1) => FP_Z(1), FP_Z(0) => FP_Z(0));
   n1 <= '0';

end SYN_pipeline;
