package myPkg is

	constant nb : integer := 14;

end myPkg;
