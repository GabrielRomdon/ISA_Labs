package my_pkg is

	constant n_levels : integer := 7;

end my_pkg;
