package CONSTANTS is
   constant NBIT_PER_BLOCK : integer :=4;
   constant NBLOCKS : integer := 16;
   constant NBIT : integer := NBLOCKS*NBIT_PER_BLOCK;
end CONSTANTS;
