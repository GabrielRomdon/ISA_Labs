package lookah_pkg is
	constant nb : integer := 14;
	constant r : integer := 7; 
	constant nb_w : integer := 15; 
	constant nb_a : integer := 14;	
	constant nb_fb : integer := 6;
end lookah_pkg;
