package myPkg is

	constant nb : integer := 14;
	constant r : integer := 3;

end myPkg;
