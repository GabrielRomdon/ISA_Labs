package lookah_pkg is
	constant nb : integer := 14;
	constant r : integer := 7; --5
	constant nb_w : integer := 15; --17vers0
	constant nb_a : integer := 14;	--22
	constant nb_fb : integer := 7;
end lookah_pkg;
