
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_FPmul is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_FPmul;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_9;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_57 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_57;

architecture SYN_BEHAVIORAL of PG_GENERAL_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_53 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_53;

architecture SYN_BEHAVIORAL of PG_GENERAL_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_49 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_49;

architecture SYN_BEHAVIORAL of PG_GENERAL_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_60 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_60;

architecture SYN_BEHAVIORAL of PG_GENERAL_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_59 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_59;

architecture SYN_BEHAVIORAL of PG_GENERAL_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_43 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_43;

architecture SYN_BEHAVIORAL of PG_GENERAL_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_44 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_44;

architecture SYN_BEHAVIORAL of PG_GENERAL_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_32 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_32;

architecture SYN_BEHAVIORAL of PG_GENERAL_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_31 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_31;

architecture SYN_BEHAVIORAL of PG_GENERAL_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_12 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_12;

architecture SYN_BEHAVIORAL of G_GENERAL_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_11 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_11;

architecture SYN_BEHAVIORAL of G_GENERAL_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_8 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_8;

architecture SYN_BEHAVIORAL of G_GENERAL_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_30 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_30;

architecture SYN_BEHAVIORAL of PG_NET_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XNOR2_X1 port map( A => A, B => n1, ZN => P_OUT);
   U3 : INV_X1 port map( A => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_50 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_50;

architecture SYN_BEHAVIORAL of PG_NET_50 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_45 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_45;

architecture SYN_BEHAVIORAL of PG_NET_45 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_42 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_42;

architecture SYN_BEHAVIORAL of PG_NET_42 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_39 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_39;

architecture SYN_BEHAVIORAL of PG_NET_39 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_38 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_38;

architecture SYN_BEHAVIORAL of PG_NET_38 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_31 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_31;

architecture SYN_BEHAVIORAL of PG_NET_31 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_25 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_25;

architecture SYN_BEHAVIORAL of PG_NET_25 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_58 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_58;

architecture SYN_BEHAVIORAL of PG_NET_58 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_57 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_57;

architecture SYN_BEHAVIORAL of PG_NET_57 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_56 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_56;

architecture SYN_BEHAVIORAL of PG_NET_56 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_55 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_55;

architecture SYN_BEHAVIORAL of PG_NET_55 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_53 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_53;

architecture SYN_BEHAVIORAL of PG_NET_53 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_52 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_52;

architecture SYN_BEHAVIORAL of PG_NET_52 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_48 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_48;

architecture SYN_BEHAVIORAL of PG_NET_48 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_47 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_47;

architecture SYN_BEHAVIORAL of PG_NET_47 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_46 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_46;

architecture SYN_BEHAVIORAL of PG_NET_46 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_41 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_41;

architecture SYN_BEHAVIORAL of PG_NET_41 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_29 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_29;

architecture SYN_BEHAVIORAL of PG_NET_29 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_24 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_24;

architecture SYN_BEHAVIORAL of PG_NET_24 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_23 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_23;

architecture SYN_BEHAVIORAL of PG_NET_23 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_21 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_21;

architecture SYN_BEHAVIORAL of PG_NET_21 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n2, ZN => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_567 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_567;

architecture SYN_BEHAVIORAL of FA_567 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_460;

architecture SYN_BEHAVIORAL of FA_460 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_477 is

   port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_477;

architecture SYN_BEHAVIORAL of FA_477 is

begin
   S_BAR <= A_BAR;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_365 is

   port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_365;

architecture SYN_BEHAVIORAL of FA_365 is

begin
   S_BAR <= A_BAR;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_577 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_577;

architecture SYN_BEHAVIORAL of FA_577 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_576 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_576;

architecture SYN_BEHAVIORAL of FA_576 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_544 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_544;

architecture SYN_BEHAVIORAL of FA_544 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_504;

architecture SYN_BEHAVIORAL of FA_504 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_481;

architecture SYN_BEHAVIORAL of FA_481 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n2, B2 => n3, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_487 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_487;

architecture SYN_BEHAVIORAL of FA_487 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_529 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_529;

architecture SYN_BEHAVIORAL of FA_529 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_505;

architecture SYN_BEHAVIORAL of FA_505 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_462;

architecture SYN_BEHAVIORAL of FA_462 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_379;

architecture SYN_BEHAVIORAL of FA_379 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n2, n3 : std_logic;

begin
   S <= S_port;
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => S_port);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_367;

architecture SYN_BEHAVIORAL of FA_367 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_542 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_542;

architecture SYN_BEHAVIORAL of FA_542 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_540 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_540;

architecture SYN_BEHAVIORAL of FA_540 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_491 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_491;

architecture SYN_BEHAVIORAL of FA_491 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_490 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_490;

architecture SYN_BEHAVIORAL of FA_490 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_489 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_489;

architecture SYN_BEHAVIORAL of FA_489 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_514 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_514;

architecture SYN_BEHAVIORAL of FA_514 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_513 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_513;

architecture SYN_BEHAVIORAL of FA_513 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_512 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_512;

architecture SYN_BEHAVIORAL of FA_512 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_510;

architecture SYN_BEHAVIORAL of FA_510 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_419;

architecture SYN_BEHAVIORAL of FA_419 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_418;

architecture SYN_BEHAVIORAL of FA_418 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_417;

architecture SYN_BEHAVIORAL of FA_417 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_416;

architecture SYN_BEHAVIORAL of FA_416 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_380;

architecture SYN_BEHAVIORAL of FA_380 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_377;

architecture SYN_BEHAVIORAL of FA_377 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_376;

architecture SYN_BEHAVIORAL of FA_376 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_375;

architecture SYN_BEHAVIORAL of FA_375 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_344;

architecture SYN_BEHAVIORAL of FA_344 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_343;

architecture SYN_BEHAVIORAL of FA_343 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_18;

architecture SYN_STRUCTURAL of RCA_generic_N4_18 is

   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102722, n_1065 : std_logic;

begin
   
   net102722 <= '0';
   FAI_1 : FA_72 port map( A => A(0), B => B(0), Ci => net102722, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_71 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_70 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_69 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1065);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_39 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_39;

architecture SYN_rtl of HA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_36 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_36;

architecture SYN_rtl of HA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_35 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_35;

architecture SYN_rtl of HA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_34 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_34;

architecture SYN_rtl of HA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_32 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_32;

architecture SYN_rtl of HA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_31 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_31;

architecture SYN_rtl of HA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_28 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_28;

architecture SYN_rtl of HA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_25 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_25;

architecture SYN_rtl of HA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_23 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_23;

architecture SYN_rtl of HA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_22 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_22;

architecture SYN_rtl of HA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_20 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_20;

architecture SYN_rtl of HA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_17 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_17;

architecture SYN_rtl of HA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_16 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_16;

architecture SYN_rtl of HA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_14 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_14;

architecture SYN_rtl of HA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_13 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_13;

architecture SYN_rtl of HA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_11 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_11;

architecture SYN_rtl of HA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_10 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_10;

architecture SYN_rtl of HA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_8 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_8;

architecture SYN_rtl of HA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_7 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_7;

architecture SYN_rtl of HA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_5 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_5;

architecture SYN_rtl of HA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_4 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_4;

architecture SYN_rtl of HA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_2 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_2;

architecture SYN_rtl of HA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_1 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_1;

architecture SYN_rtl of HA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_536 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_536;

architecture SYN_BEHAVIORAL of FA_536 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_56 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_56;

architecture SYN_BEHAVIORAL of PG_GENERAL_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_32 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_32;

architecture SYN_BEHAVIORAL of PG_NET_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_28 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_28;

architecture SYN_BEHAVIORAL of PG_NET_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_26 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_26;

architecture SYN_BEHAVIORAL of PG_NET_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_341;

architecture SYN_BEHAVIORAL of FA_341 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);
   U7 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);
   U2 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U4 : INV_X1 port map( A => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_43 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co_BAR : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => Co_BAR);
   U6 : XOR2_X1 port map( A => n4, B => B, Z => S);
   U1 : INV_X1 port map( A => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U7 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n6, n8, n9, n10 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n6, ZN => Co);
   U6 : NAND2_X1 port map( A1 => n8, A2 => B, ZN => n6);
   U8 : INV_X1 port map( A => n2, ZN => n8);
   U9 : NAND2_X1 port map( A1 => Ci, A2 => n10, ZN => n9);
   U10 : INV_X1 port map( A => n4, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);
   U3 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U4 : INV_X1 port map( A => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n7, Z => S);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n7, n9, n10, n12 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U7 : XOR2_X1 port map( A => Ci, B => n12, Z => S);
   U3 : NAND2_X1 port map( A1 => n10, A2 => n7, ZN => Co);
   U5 : NAND2_X1 port map( A1 => n9, A2 => B, ZN => n7);
   U9 : INV_X1 port map( A => n2, ZN => n9);
   U10 : NAND2_X1 port map( A1 => Ci, A2 => n12, ZN => n10);
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n3);
   U3 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n3, B2 => n2, ZN => Co);
   U7 : INV_X1 port map( A => n5, ZN => n6);
   U8 : XOR2_X1 port map( A => Ci, B => n6, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_port, n2, n3 : std_logic;

begin
   S <= S_port;
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => S_port);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => S_port, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   U6 : INV_X1 port map( A => n4, ZN => n5);
   U7 : XOR2_X1 port map( A => Ci, B => n5, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n5, ZN => Co);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U2 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U3 : INV_X1 port map( A => Ci, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U2 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  clk : in std_logic);

end MUX21_GENERIC_N4_5;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_5 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal n29, n30, n31, n32, n33, n_1091, n_1092, n_1093, n_1094, n_1095 : 
      std_logic;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => n30, B => n32, S => n29, Z => Y(0));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => n31, B => n33, S => n29, Z => Y(2));
   MY_CLK_r_REG351_S3 : DFF_X1 port map( D => A(2), CK => clk, Q => n33, QN => 
                           n_1091);
   MY_CLK_r_REG352_S3 : DFF_X1 port map( D => A(0), CK => clk, Q => n32, QN => 
                           n_1092);
   MY_CLK_r_REG350_S3 : DFF_X1 port map( D => B(2), CK => clk, Q => n31, QN => 
                           n_1093);
   MY_CLK_r_REG349_S3 : DFF_X1 port map( D => B(0), CK => clk, Q => n30, QN => 
                           n_1094);
   MY_CLK_r_REG248_S3 : DFF_X1 port map( D => SEL, CK => clk, Q => n29, QN => 
                           n_1095);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_9;

architecture SYN_STRUCTURAL of RCA_generic_N4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102723, n_1098 : std_logic;

begin
   
   net102723 <= '0';
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => net102723, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1098);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_10;

architecture SYN_STRUCTURAL of RCA_generic_N4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102721, n_1101 : std_logic;

begin
   
   net102721 <= '0';
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => net102721, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1101);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  clk : in std_logic);

end MUX21_GENERIC_N4_6;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_11;

architecture SYN_STRUCTURAL of RCA_generic_N4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102724, n_1104 : std_logic;

begin
   
   net102724 <= '0';
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => net102724, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), S => S(1), Co => CTMP_2_port, 
                           Ci_BAR => CTMP_1_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1104);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_12;

architecture SYN_STRUCTURAL of RCA_generic_N4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102721, n_1107 : std_logic;

begin
   
   net102721 <= '0';
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => net102721, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1107);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0);  clk : in std_logic);

end MUX21_GENERIC_N4_7;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_13;

architecture SYN_STRUCTURAL of RCA_generic_N4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102726, n_1110 : std_logic;

begin
   
   net102726 <= '0';
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => net102726, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1110);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_14;

architecture SYN_STRUCTURAL of RCA_generic_N4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102720, n_1113 : std_logic;

begin
   
   net102720 <= '0';
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => net102720, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1113);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_8;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_15;

architecture SYN_STRUCTURAL of RCA_generic_N4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102727, n_1116 : std_logic;

begin
   
   net102727 <= '0';
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => net102727, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1116);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_16;

architecture SYN_STRUCTURAL of RCA_generic_N4_16 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102720, n_1119 : std_logic;

begin
   
   net102720 <= '0';
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => net102720, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1119);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_17;

architecture SYN_STRUCTURAL of RCA_generic_N4_17 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102729, n_1122 : std_logic;

begin
   
   net102729 <= '0';
   FAI_1 : FA_68 port map( A => A(0), B => B(0), Ci => net102729, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_67 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_66 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_65 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1122);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_10;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));
   U2 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_19;

architecture SYN_STRUCTURAL of RCA_generic_N4_19 is

   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102730, n_1125 : std_logic;

begin
   
   net102730 <= '0';
   FAI_1 : FA_76 port map( A => A(0), B => B(0), Ci => net102730, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_75 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_74 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_73 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1125);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_20;

architecture SYN_STRUCTURAL of RCA_generic_N4_20 is

   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102722, n_1128 : std_logic;

begin
   
   net102722 <= '0';
   FAI_1 : FA_80 port map( A => A(0), B => B(0), Ci => net102722, S => S(0), Co
                           => CTMP_1_port);
   FAI_2 : FA_79 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_78 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_77 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1128);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MUX21_GENERIC_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_N4_11;

architecture SYN_BEHAVIORAL of MUX21_GENERIC_N4_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U3 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_21;

architecture SYN_STRUCTURAL of RCA_generic_N4_21 is

   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102732, n_1139, n_1140, 
      n_1141 : std_logic;

begin
   
   net102732 <= '0';
   FAI_1 : FA_84 port map( A => A(0), B => B(0), Ci => net102732, S => n_1139, 
                           Co => CTMP_1_port);
   FAI_2 : FA_83 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => n_1140
                           , Co => CTMP_2_port);
   FAI_3 : FA_82 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_81 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1141);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity RCA_generic_N4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_generic_N4_22;

architecture SYN_STRUCTURAL of RCA_generic_N4_22 is

   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port, net102733, n_1146, n_1147, 
      n_1148 : std_logic;

begin
   
   net102733 <= '0';
   FAI_1 : FA_88 port map( A => A(0), B => B(0), Ci => net102733, S => n_1146, 
                           Co => CTMP_1_port);
   FAI_2 : FA_87 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => n_1147
                           , Co => CTMP_2_port);
   FAI_3 : FA_86 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_85 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => n_1148);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  clk : in std_logic);

end carry_select_N4_5;

architecture SYN_STRUCTURAL of carry_select_N4_5 is

   component MUX21_GENERIC_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  clk : in std_logic);
   end component;
   
   component RCA_generic_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n10, n11, n12, n13
      , n14, n15, n16, n17, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, 
      n_1155, n_1156, n_1157, n_1158 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   MY_CLK_r_REG366_S2 : DFF_X1 port map( D => A(3), CK => clk, Q => n17, QN => 
                           n_1149);
   MY_CLK_r_REG367_S2 : DFF_X1 port map( D => A(2), CK => clk, Q => n16, QN => 
                           n_1150);
   MY_CLK_r_REG359_S2 : DFF_X1 port map( D => A(1), CK => clk, Q => n15, QN => 
                           n_1151);
   MY_CLK_r_REG360_S2 : DFF_X1 port map( D => A(0), CK => clk, Q => n14, QN => 
                           n_1152);
   MY_CLK_r_REG368_S2 : DFF_X1 port map( D => B(3), CK => clk, Q => n13, QN => 
                           n_1153);
   MY_CLK_r_REG358_S2 : DFF_X1 port map( D => B(2), CK => clk, Q => n12, QN => 
                           n_1154);
   MY_CLK_r_REG361_S2 : DFF_X1 port map( D => B(1), CK => clk, Q => n11, QN => 
                           n_1155);
   MY_CLK_r_REG348_S2 : DFF_X1 port map( D => B(0), CK => clk, Q => n10, QN => 
                           n_1156);
   ADDER0 : RCA_generic_N4_10 port map( A(3) => n17, A(2) => n16, A(1) => n15, 
                           A(0) => n14, B(3) => n13, B(2) => n12, B(1) => n11, 
                           B(0) => n10, Ci => X_Logic0_port, S(3) => S0_3_port,
                           S(2) => S0_2_port, S(1) => S0_1_port, S(0) => 
                           S0_0_port, Co => n_1157);
   ADDER1 : RCA_generic_N4_9 port map( A(3) => n17, A(2) => n16, A(1) => n15, 
                           A(0) => n14, B(3) => n13, B(2) => n12, B(1) => n11, 
                           B(0) => n10, Ci => X_Logic1_port, S(3) => S1_3_port,
                           S(2) => S1_2_port, S(1) => S1_1_port, S(0) => 
                           S1_0_port, Co => n_1158);
   MUX : MUX21_GENERIC_N4_5 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0), clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  clk : in std_logic);

end carry_select_N4_6;

architecture SYN_STRUCTURAL of carry_select_N4_6 is

   component MUX21_GENERIC_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  clk : in std_logic);
   end component;
   
   component RCA_generic_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1159, n_1160 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1159);
   ADDER1 : RCA_generic_N4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1160);
   MUX : MUX21_GENERIC_N4_6 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0), clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  clk : in std_logic);

end carry_select_N4_7;

architecture SYN_STRUCTURAL of carry_select_N4_7 is

   component MUX21_GENERIC_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0);  clk : in std_logic);
   end component;
   
   component RCA_generic_N4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1161, n_1162 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1161);
   ADDER1 : RCA_generic_N4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1162);
   MUX : MUX21_GENERIC_N4_7 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0), clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_8;

architecture SYN_STRUCTURAL of carry_select_N4_8 is

   component MUX21_GENERIC_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1163, n_1164 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1163);
   ADDER1 : RCA_generic_N4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1164);
   MUX : MUX21_GENERIC_N4_8 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_9;

architecture SYN_STRUCTURAL of carry_select_N4_9 is

   component MUX21_GENERIC_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1165, n_1166 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1165);
   ADDER1 : RCA_generic_N4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1166);
   MUX : MUX21_GENERIC_N4_9 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_10;

architecture SYN_STRUCTURAL of carry_select_N4_10 is

   component MUX21_GENERIC_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, n_1167, n_1168 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ADDER0 : RCA_generic_N4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => n_1167);
   ADDER1 : RCA_generic_N4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => n_1168);
   MUX : MUX21_GENERIC_N4_10 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => S1_1_port, A(0) => S1_0_port, B(3) => 
                           S0_3_port, B(2) => S0_2_port, B(1) => S0_1_port, 
                           B(0) => S0_0_port, SEL => Ci, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity carry_select_N4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0));

end carry_select_N4_11;

architecture SYN_STRUCTURAL of carry_select_N4_11 is

   component MUX21_GENERIC_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_generic_N4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, S0_3_port, S0_2_port, S1_3_port, 
      S1_2_port, n1, n2, n3, n4, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176
      , n_1177, n_1178 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n1 <= '0';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   ADDER0 : RCA_generic_N4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => n_1171, S(0) 
                           => n_1172, Co => n_1173);
   ADDER1 : RCA_generic_N4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => n_1174, S(0) 
                           => n_1175, Co => n_1176);
   MUX : MUX21_GENERIC_N4_11 port map( A(3) => S1_3_port, A(2) => S1_2_port, 
                           A(1) => n1, A(0) => n2, B(3) => S0_3_port, B(2) => 
                           S0_2_port, B(1) => n3, B(0) => n4, SEL => Ci, Y(3) 
                           => S(3), Y(2) => S(2), Y(1) => n_1177, Y(0) => 
                           n_1178);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_6 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_6;

architecture SYN_BEHAVIORAL of G_GENERAL_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => G_k_1j, A2 => PG_ik(0), ZN => n2);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => G_ij);
   U3 : INV_X1 port map( A => PG_ik(1), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_7 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_7;

architecture SYN_BEHAVIORAL of G_GENERAL_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => G_ij);
   U2 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_9 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_9;

architecture SYN_BEHAVIORAL of G_GENERAL_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : OR2_X2 port map( A1 => PG_ik(1), A2 => n1, ZN => G_ij);
   U2 : AND2_X1 port map( A1 => PG_ik(0), A2 => G_k_1j, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_10 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_10;

architecture SYN_BEHAVIORAL of G_GENERAL_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => PG_ik(1), A2 => n5, ZN => G_ij);
   U2 : AND2_X1 port map( A1 => PG_ik(0), A2 => G_k_1j, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_8 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_8;

architecture SYN_BEHAVIORAL of PG_GENERAL_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U1 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => PG_ij(1));
   U2 : INV_X1 port map( A => PG_ik(1), ZN => n2);
   U4 : NAND2_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(0), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_9 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_9;

architecture SYN_BEHAVIORAL of PG_GENERAL_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U1 : NAND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n2);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => PG_ij(1));
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_10 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_10;

architecture SYN_BEHAVIORAL of PG_GENERAL_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_13 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic;  clk : in std_logic);

end G_GENERAL_13;

architecture SYN_BEHAVIORAL of G_GENERAL_13 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n_1179 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n3, B2 => PG_ik(0), A => PG_ik(1), ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);
   MY_CLK_r_REG570_S2 : DFF_X1 port map( D => G_k_1j, CK => clk, Q => n3, QN =>
                           n_1179);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_14 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_14;

architecture SYN_BEHAVIORAL of PG_GENERAL_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U1 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => PG_ij(1));
   U2 : NAND2_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(0), ZN => n2);
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_15 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_15;

architecture SYN_BEHAVIORAL of PG_GENERAL_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : NAND2_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(0), ZN => n3);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => PG_ij(1));
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_16 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_16;

architecture SYN_BEHAVIORAL of PG_GENERAL_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U3 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U1 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => PG_ij(1));
   U2 : NAND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n3);
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_17 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_17;

architecture SYN_BEHAVIORAL of PG_GENERAL_17 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n_1180, n_1181 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n4, A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AND2_X1 port map( A1 => n5, A2 => PG_ik(0), ZN => n3);
   U3 : OR2_X1 port map( A1 => PG_ik(1), A2 => n3, ZN => PG_ij(1));
   MY_CLK_r_REG536_S2 : DFF_X1 port map( D => PG_k_1j(1), CK => clk, Q => n5, 
                           QN => n_1180);
   MY_CLK_r_REG537_S2 : DFF_X1 port map( D => PG_k_1j(0), CK => clk, Q => n4, 
                           QN => n_1181);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_15 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_15;

architecture SYN_BEHAVIORAL of G_GENERAL_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => G_k_1j, B2 => PG_ik(0), A => PG_ik(1), ZN => 
                           n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_23 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_23;

architecture SYN_BEHAVIORAL of PG_GENERAL_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_24 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_24;

architecture SYN_BEHAVIORAL of PG_GENERAL_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U1 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => PG_ij(1));
   U2 : INV_X1 port map( A => PG_ik(1), ZN => n2);
   U4 : NAND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_25 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_25;

architecture SYN_BEHAVIORAL of PG_GENERAL_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => PG_ij(1));
   U3 : INV_X1 port map( A => PG_ik(1), ZN => n3);
   U4 : NAND2_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(0), ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_26 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_26;

architecture SYN_BEHAVIORAL of PG_GENERAL_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net39840, n1, n2 : std_logic;

begin
   
   U2 : OAI21_X1 port map( B1 => n1, B2 => net39840, A => n2, ZN => PG_ij(1));
   U3 : INV_X1 port map( A => PG_k_1j(1), ZN => n1);
   U4 : INV_X1 port map( A => PG_ik(0), ZN => net39840);
   U5 : INV_X1 port map( A => PG_ik(1), ZN => n2);
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_27 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_27;

architecture SYN_BEHAVIORAL of PG_GENERAL_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6 : std_logic;

begin
   
   U5 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U1 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => PG_ij(1));
   U2 : NAND2_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(0), ZN => n5);
   U3 : INV_X1 port map( A => PG_ik(1), ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_28 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_28;

architecture SYN_BEHAVIORAL of PG_GENERAL_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U1 : INV_X1 port map( A => PG_ik(1), ZN => n4);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => PG_ij(1));
   U4 : NAND2_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(0), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_29 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_29;

architecture SYN_BEHAVIORAL of PG_GENERAL_29 is

   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7, n_1182, n_1183, n_1184 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n5, A2 => n7, ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => n6, B2 => n7, A => PG_ik(1), ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));
   MY_CLK_r_REG473_S2 : DFF_X1 port map( D => PG_k_1j(1), CK => clk, Q => n6, 
                           QN => n_1182);
   MY_CLK_r_REG474_S2 : DFF_X1 port map( D => PG_k_1j(0), CK => clk, Q => n5, 
                           QN => n_1183);
   MY_CLK_r_REG461_S2 : DFF_X2 port map( D => PG_ik(0), CK => clk, Q => n7, QN 
                           => n_1184);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_30 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_30;

architecture SYN_BEHAVIORAL of PG_GENERAL_30 is

   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6, n7, n8, n9, n_1185, n_1186, n_1187, n_1188 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n6, A2 => n8, ZN => PG_ij(0));
   U2 : OR2_X1 port map( A1 => n4, A2 => n9, ZN => PG_ij(1));
   U3 : AND2_X1 port map( A1 => n7, A2 => n8, ZN => n4);
   MY_CLK_r_REG501_S2 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n8, QN 
                           => n_1185);
   MY_CLK_r_REG514_S2 : DFF_X1 port map( D => PG_k_1j(1), CK => clk, Q => n7, 
                           QN => n_1186);
   MY_CLK_r_REG515_S2 : DFF_X1 port map( D => PG_k_1j(0), CK => clk, Q => n6, 
                           QN => n_1187);
   MY_CLK_r_REG500_S2 : DFF_X2 port map( D => PG_ik(1), CK => clk, Q => n9, QN 
                           => n_1188);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_16 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic;  clk : in std_logic);

end G_GENERAL_16;

architecture SYN_BEHAVIORAL of G_GENERAL_16 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n7, n_1189, n_1190, n_1191 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n5, B2 => n6, A => n7, ZN => n1);
   U2 : INV_X1 port map( A => n1, ZN => G_ij);
   MY_CLK_r_REG616_S1 : DFF_X1 port map( D => PG_ik(1), CK => clk, Q => n7, QN 
                           => n_1189);
   MY_CLK_r_REG617_S1 : DFF_X1 port map( D => PG_ik(0), CK => clk, Q => n6, QN 
                           => n_1190);
   MY_CLK_r_REG634_S1 : DFF_X1 port map( D => G_k_1j, CK => clk, Q => n5, QN =>
                           n_1191);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_45 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_45;

architecture SYN_BEHAVIORAL of PG_GENERAL_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PG_ij(1));
   U2 : INV_X1 port map( A => PG_ik(0), ZN => n1);
   U3 : INV_X1 port map( A => PG_k_1j(1), ZN => n2);
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n3);
   U5 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_46 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_46;

architecture SYN_BEHAVIORAL of PG_GENERAL_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => PG_ij(1));
   U2 : INV_X1 port map( A => PG_ik(0), ZN => n1);
   U3 : INV_X1 port map( A => PG_k_1j(1), ZN => n2);
   U4 : INV_X1 port map( A => PG_ik(1), ZN => n3);
   U6 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_47 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_47;

architecture SYN_BEHAVIORAL of PG_GENERAL_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : INV_X1 port map( A => PG_ik(1), ZN => n3);
   U3 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => PG_ij(1));
   U4 : NAND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_48 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_48;

architecture SYN_BEHAVIORAL of PG_GENERAL_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U3 : OAI22_X1 port map( A1 => PG_k_1j(1), A2 => PG_ik(1), B1 => PG_ik(0), B2
                           => PG_ik(1), ZN => n2);
   U4 : INV_X1 port map( A => n2, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_50 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_50;

architecture SYN_BEHAVIORAL of PG_GENERAL_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net39810, n1, n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : OAI21_X1 port map( B1 => net39810, B2 => n1, A => n2, ZN => PG_ij(1));
   U3 : INV_X1 port map( A => PG_ik(0), ZN => net39810);
   U4 : INV_X1 port map( A => PG_k_1j(1), ZN => n1);
   U5 : INV_X1 port map( A => PG_ik(1), ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_51 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_51;

architecture SYN_BEHAVIORAL of PG_GENERAL_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => PG_ij(1));
   U4 : NAND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n4);
   U3 : INV_X1 port map( A => PG_ik(1), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_52 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_52;

architecture SYN_BEHAVIORAL of PG_GENERAL_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U1 : INV_X1 port map( A => PG_ik(1), ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => PG_ij(1));
   U4 : NAND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(1), ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_54 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_54;

architecture SYN_BEHAVIORAL of PG_GENERAL_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : OAI22_X1 port map( A1 => PG_ik(0), A2 => PG_ik(1), B1 => PG_k_1j(1), B2
                           => PG_ik(1), ZN => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_55 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0);  clk : in std_logic);

end PG_GENERAL_55;

architecture SYN_BEHAVIORAL of PG_GENERAL_55 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n_1192 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   MY_CLK_r_REG460_S2 : DFF_X1 port map( D => n1, CK => clk, Q => n_1192, QN =>
                           PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_58 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_58;

architecture SYN_BEHAVIORAL of PG_GENERAL_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_ik(0), A2 => PG_k_1j(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_61 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_61;

architecture SYN_BEHAVIORAL of PG_GENERAL_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_ik(0), B2 => PG_k_1j(1), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_62 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_62;

architecture SYN_BEHAVIORAL of PG_GENERAL_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_GENERAL_0 is

   port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
         std_logic_vector (1 downto 0));

end PG_GENERAL_0;

architecture SYN_BEHAVIORAL of PG_GENERAL_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => PG_k_1j(0), A2 => PG_ik(0), ZN => PG_ij(0));
   U2 : AOI21_X1 port map( B1 => PG_k_1j(1), B2 => PG_ik(0), A => PG_ik(1), ZN 
                           => n1);
   U3 : INV_X1 port map( A => n1, ZN => PG_ij(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity G_GENERAL_0 is

   port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
         G_ij : out std_logic);

end G_GENERAL_0;

architecture SYN_BEHAVIORAL of G_GENERAL_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => G_k_1j, A2 => PG_ik(0), ZN => G_ij);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_22 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_22;

architecture SYN_BEHAVIORAL of PG_NET_22 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n2, ZN => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_27 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_27;

architecture SYN_BEHAVIORAL of PG_NET_27 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net27166, net27167 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => net27166);
   U3 : INV_X1 port map( A => B, ZN => net27167);
   U4 : NOR2_X1 port map( A1 => net27166, A2 => net27167, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_33 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_33;

architecture SYN_BEHAVIORAL of PG_NET_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U3 : XNOR2_X1 port map( A => n2, B => A, ZN => P_OUT);
   U4 : INV_X1 port map( A => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_34 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_34;

architecture SYN_BEHAVIORAL of PG_NET_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U3 : XNOR2_X1 port map( A => n2, B => A, ZN => P_OUT);
   U4 : INV_X1 port map( A => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_35 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_35;

architecture SYN_BEHAVIORAL of PG_NET_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net27183, n1 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U3 : INV_X1 port map( A => B, ZN => net27183);
   U4 : NOR2_X1 port map( A1 => n1, A2 => net27183, ZN => G_OUT);
   U5 : INV_X1 port map( A => A, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_36 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_36;

architecture SYN_BEHAVIORAL of PG_NET_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_37 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_37;

architecture SYN_BEHAVIORAL of PG_NET_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U3 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_40 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_40;

architecture SYN_BEHAVIORAL of PG_NET_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_43 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_43;

architecture SYN_BEHAVIORAL of PG_NET_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_44 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_44;

architecture SYN_BEHAVIORAL of PG_NET_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_49 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_49;

architecture SYN_BEHAVIORAL of PG_NET_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => G_OUT);
   U1 : XNOR2_X1 port map( A => n3, B => A, ZN => P_OUT);
   U3 : INV_X1 port map( A => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_51 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_51;

architecture SYN_BEHAVIORAL of PG_NET_51 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => P_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_54 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_54;

architecture SYN_BEHAVIORAL of PG_NET_54 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_59 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
         std_logic);

end PG_NET_59;

architecture SYN_BEHAVIORAL of PG_NET_59 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n_1194 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => n2, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => n2, B => A, Z => P_OUT);
   MY_CLK_r_REG604_S1 : DFF_X1 port map( D => B, CK => clk, Q => n2, QN => 
                           n_1194);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_60 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
         std_logic);

end PG_NET_60;

architecture SYN_BEHAVIORAL of PG_NET_60 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n_1195 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => n2, ZN => G_OUT);
   U2 : XOR2_X1 port map( A => n2, B => A, Z => P_OUT);
   MY_CLK_r_REG618_S1 : DFF_X1 port map( D => B, CK => clk, Q => n2, QN => 
                           n_1195);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_61 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_61;

architecture SYN_BEHAVIORAL of PG_NET_61 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_62 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_62;

architecture SYN_BEHAVIORAL of PG_NET_62 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P_OUT);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_63 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_63;

architecture SYN_BEHAVIORAL of PG_NET_63 is

begin
   P_OUT <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PG_NET_0 is

   port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);

end PG_NET_0;

architecture SYN_BEHAVIORAL of PG_NET_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n2);
   U3 : INV_X1 port map( A => B, ZN => n1);
   U4 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => G_OUT);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic_vector 
         (15 downto 0);  S : out std_logic_vector (63 downto 0);  clk : in 
         std_logic);

end SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16;

architecture SYN_STRUCTURAL of SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16 is

   component carry_select_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  clk : in std_logic);
   end component;
   
   component carry_select_N4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   signal n_1318, n_1319 : std_logic;

begin
   
   CS_5 : carry_select_N4_11 port map( A(3) => A(23), A(2) => A(22), A(1) => 
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Ci => Ci(5), S(3) => 
                           S(23), S(2) => S(22), S(1) => n_1318, S(0) => n_1319
                           );
   CS_6 : carry_select_N4_10 port map( A(3) => A(27), A(2) => A(26), A(1) => 
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Ci => Ci(6), S(3) => 
                           S(27), S(2) => S(26), S(1) => S(25), S(0) => S(24));
   CS_7 : carry_select_N4_9 port map( A(3) => A(31), A(2) => A(30), A(1) => 
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Ci => Ci(7), S(3) => 
                           S(31), S(2) => S(30), S(1) => S(29), S(0) => S(28));
   CS_8 : carry_select_N4_8 port map( A(3) => A(35), A(2) => A(34), A(1) => 
                           A(33), A(0) => A(32), B(3) => B(35), B(2) => B(34), 
                           B(1) => B(33), B(0) => B(32), Ci => Ci(8), S(3) => 
                           S(35), S(2) => S(34), S(1) => S(33), S(0) => S(32));
   CS_9 : carry_select_N4_7 port map( A(3) => A(39), A(2) => A(38), A(1) => 
                           A(37), A(0) => A(36), B(3) => B(39), B(2) => B(38), 
                           B(1) => B(37), B(0) => B(36), Ci => Ci(9), S(3) => 
                           S(39), S(2) => S(38), S(1) => S(37), S(0) => S(36), 
                           clk => clk);
   CS_10 : carry_select_N4_6 port map( A(3) => A(43), A(2) => A(42), A(1) => 
                           A(41), A(0) => A(40), B(3) => B(43), B(2) => B(42), 
                           B(1) => B(41), B(0) => B(40), Ci => Ci(10), S(3) => 
                           S(43), S(2) => S(42), S(1) => S(41), S(0) => S(40), 
                           clk => clk);
   CS_11 : carry_select_N4_5 port map( A(3) => A(47), A(2) => A(46), A(1) => 
                           A(45), A(0) => A(44), B(3) => B(47), B(2) => B(46), 
                           B(1) => B(45), B(0) => B(44), Ci => Ci(11), S(3) => 
                           S(47), S(2) => S(46), S(1) => S(45), S(0) => S(44), 
                           clk => clk);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (16 downto 0);  clk : in std_logic);

end CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4;

architecture SYN_STRUCTURAL of CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component G_GENERAL_6
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_7
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_8
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_9
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_10
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_11
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component G_GENERAL_12
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_8
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_9
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_10
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_13
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic;  clk : in std_logic);
   end component;
   
   component PG_GENERAL_14
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_15
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_16
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_17
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component G_GENERAL_15
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_GENERAL_23
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_24
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_25
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_26
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_27
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_28
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_29
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_30
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_31
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_32
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_16
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic;  clk : in std_logic);
   end component;
   
   component PG_GENERAL_43
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_44
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_45
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_46
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_47
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_48
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_49
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_50
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_51
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_52
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_53
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_54
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_55
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0);  clk : in std_logic);
   end component;
   
   component PG_GENERAL_56
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_57
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_58
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_59
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_60
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_61
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_62
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component PG_GENERAL_0
      port( PG_ik, PG_k_1j : in std_logic_vector (1 downto 0);  PG_ij : out 
            std_logic_vector (1 downto 0));
   end component;
   
   component G_GENERAL_0
      port( PG_ik : in std_logic_vector (1 downto 0);  G_k_1j : in std_logic;  
            G_ij : out std_logic);
   end component;
   
   component PG_NET_21
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_22
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_23
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_24
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_25
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_26
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_27
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_28
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_29
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_30
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_31
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_32
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_33
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_34
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_35
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_36
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_37
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_38
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_39
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_40
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_41
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_42
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_43
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_44
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_45
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_46
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_47
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_48
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_49
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_50
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_51
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_52
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_53
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_54
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_55
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_56
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_57
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_58
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_59
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component PG_NET_60
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component PG_NET_61
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_62
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_63
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component PG_NET_0
      port( A, B : in std_logic;  G_OUT, P_OUT : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n8, n9, n10, n11, lev_i_out_4_44_1_port, lev_i_out_4_44_0_port, 
      lev_i_out_4_32_1_port, lev_i_out_4_32_0_port, lev_i_out_4_28_1_port, 
      lev_i_out_4_28_0_port, lev_i_out_3_40_1_port, lev_i_out_3_40_0_port, 
      lev_i_out_3_32_1_port, lev_i_out_3_32_0_port, lev_i_out_3_24_1_port, 
      lev_i_out_3_24_0_port, lev_i_out_3_16_1_port, lev_i_out_3_16_0_port, 
      lev_i_out_2_44_1_port, lev_i_out_2_44_0_port, lev_i_out_2_40_1_port, 
      lev_i_out_2_40_0_port, lev_i_out_2_36_1_port, lev_i_out_2_36_0_port, 
      lev_i_out_2_32_1_port, lev_i_out_2_32_0_port, lev_i_out_2_28_0_port, 
      lev_i_out_2_24_1_port, lev_i_out_2_24_0_port, lev_i_out_2_20_1_port, 
      lev_i_out_2_20_0_port, lev_i_out_2_16_1_port, lev_i_out_2_16_0_port, 
      lev_i_out_2_12_1_port, lev_i_out_2_12_0_port, lev_i_out_2_8_1_port, 
      lev_i_out_2_8_0_port, lev_i_out_1_44_1_port, lev_i_out_1_44_0_port, 
      lev_i_out_1_42_1_port, lev_i_out_1_42_0_port, lev_i_out_1_40_1_port, 
      lev_i_out_1_40_0_port, lev_i_out_1_38_1_port, lev_i_out_1_38_0_port, 
      lev_i_out_1_36_1_port, lev_i_out_1_36_0_port, lev_i_out_1_34_1_port, 
      lev_i_out_1_34_0_port, lev_i_out_1_32_1_port, lev_i_out_1_32_0_port, 
      lev_i_out_1_30_1_port, lev_i_out_1_30_0_port, lev_i_out_1_28_1_port, 
      lev_i_out_1_28_0_port, lev_i_out_1_26_1_port, lev_i_out_1_26_0_port, 
      lev_i_out_1_24_1_port, lev_i_out_1_24_0_port, lev_i_out_1_22_1_port, 
      lev_i_out_1_22_0_port, lev_i_out_1_20_1_port, lev_i_out_1_20_0_port, 
      lev_i_out_1_18_1_port, lev_i_out_1_18_0_port, lev_i_out_1_16_1_port, 
      lev_i_out_1_16_0_port, lev_i_out_1_14_1_port, lev_i_out_1_14_0_port, 
      lev_i_out_1_12_1_port, lev_i_out_1_12_0_port, lev_i_out_1_10_1_port, 
      lev_i_out_1_10_0_port, lev_i_out_1_8_1_port, lev_i_out_1_8_0_port, 
      lev_i_out_1_6_1_port, lev_i_out_1_6_0_port, lev_i_out_1_4_1_port, 
      lev_i_out_1_4_0_port, lev_i_out_1_2_1_port, lev_i_out_0_44_1_port, 
      lev_i_out_0_44_0_port, lev_i_out_0_43_1_port, lev_i_out_0_43_0_port, 
      lev_i_out_0_42_1_port, lev_i_out_0_42_0_port, lev_i_out_0_41_1_port, 
      lev_i_out_0_41_0_port, lev_i_out_0_40_1_port, lev_i_out_0_40_0_port, 
      lev_i_out_0_39_1_port, lev_i_out_0_39_0_port, lev_i_out_0_38_1_port, 
      lev_i_out_0_38_0_port, lev_i_out_0_37_1_port, lev_i_out_0_37_0_port, 
      lev_i_out_0_36_1_port, lev_i_out_0_36_0_port, lev_i_out_0_35_1_port, 
      lev_i_out_0_35_0_port, lev_i_out_0_34_1_port, lev_i_out_0_34_0_port, 
      lev_i_out_0_33_1_port, lev_i_out_0_33_0_port, lev_i_out_0_32_1_port, 
      lev_i_out_0_32_0_port, lev_i_out_0_31_1_port, lev_i_out_0_31_0_port, 
      lev_i_out_0_30_1_port, lev_i_out_0_30_0_port, lev_i_out_0_29_1_port, 
      lev_i_out_0_29_0_port, lev_i_out_0_28_1_port, lev_i_out_0_28_0_port, 
      lev_i_out_0_27_1_port, lev_i_out_0_27_0_port, lev_i_out_0_26_1_port, 
      lev_i_out_0_26_0_port, lev_i_out_0_25_1_port, lev_i_out_0_25_0_port, 
      lev_i_out_0_24_1_port, lev_i_out_0_24_0_port, lev_i_out_0_23_1_port, 
      lev_i_out_0_23_0_port, lev_i_out_0_22_1_port, lev_i_out_0_22_0_port, 
      lev_i_out_0_21_1_port, lev_i_out_0_21_0_port, lev_i_out_0_20_1_port, 
      lev_i_out_0_20_0_port, lev_i_out_0_19_1_port, lev_i_out_0_19_0_port, 
      lev_i_out_0_18_1_port, lev_i_out_0_18_0_port, lev_i_out_0_17_1_port, 
      lev_i_out_0_17_0_port, lev_i_out_0_16_1_port, lev_i_out_0_16_0_port, 
      lev_i_out_0_15_1_port, lev_i_out_0_15_0_port, lev_i_out_0_14_1_port, 
      lev_i_out_0_14_0_port, lev_i_out_0_13_1_port, lev_i_out_0_13_0_port, 
      lev_i_out_0_12_1_port, lev_i_out_0_12_0_port, lev_i_out_0_11_1_port, 
      lev_i_out_0_11_0_port, lev_i_out_0_10_1_port, lev_i_out_0_10_0_port, 
      lev_i_out_0_9_1_port, lev_i_out_0_9_0_port, lev_i_out_0_8_1_port, 
      lev_i_out_0_8_0_port, lev_i_out_0_7_1_port, lev_i_out_0_7_0_port, 
      lev_i_out_0_6_1_port, lev_i_out_0_6_0_port, lev_i_out_0_5_1_port, 
      lev_i_out_0_5_0_port, lev_i_out_0_4_1_port, lev_i_out_0_4_0_port, 
      lev_i_out_0_3_1_port, lev_i_out_0_3_0_port, lev_i_out_0_2_0_port, 
      lev_i_out_0_1_1_port, net102734, net102735, n14, n15, n3, n_1372, n_1373 
      : std_logic;

begin
   Co <= ( Co(16), Co(15), Co(14), Co(13), Co(12), Co(11), Co(10), Co(9), Co(8)
      , Co(7), Co(6), Co(5), Co(4), Co(3), Co(2), Co(1), Co(0) );
   
   net102734 <= '0';
   net102735 <= '0';
   U4 : CLKBUF_X1 port map( A => lev_i_out_2_28_0_port, Z => n15);
   U1 : BUF_X1 port map( A => lev_i_out_3_24_1_port, Z => n14);
   PG_NETWORK_0_1 : PG_NET_0 port map( A => A(0), B => B(0), G_OUT => 
                           lev_i_out_0_1_1_port, P_OUT => n_1372);
   PG_NETWORK_0_2 : PG_NET_63 port map( A => A(1), B => net102735, G_OUT => 
                           n_1373, P_OUT => lev_i_out_0_2_0_port);
   PG_NETWORK_0_3 : PG_NET_62 port map( A => A(2), B => B(2), G_OUT => 
                           lev_i_out_0_3_1_port, P_OUT => lev_i_out_0_3_0_port)
                           ;
   PG_NETWORK_0_4 : PG_NET_61 port map( A => A(3), B => B(3), G_OUT => 
                           lev_i_out_0_4_1_port, P_OUT => lev_i_out_0_4_0_port)
                           ;
   PG_NETWORK_0_5 : PG_NET_60 port map( A => A(4), B => B(4), G_OUT => 
                           lev_i_out_0_5_1_port, P_OUT => lev_i_out_0_5_0_port,
                           clk => clk);
   PG_NETWORK_0_6 : PG_NET_59 port map( A => A(5), B => B(5), G_OUT => 
                           lev_i_out_0_6_1_port, P_OUT => lev_i_out_0_6_0_port,
                           clk => clk);
   PG_NETWORK_0_7 : PG_NET_58 port map( A => A(6), B => B(6), G_OUT => 
                           lev_i_out_0_7_1_port, P_OUT => lev_i_out_0_7_0_port)
                           ;
   PG_NETWORK_0_8 : PG_NET_57 port map( A => A(7), B => B(7), G_OUT => 
                           lev_i_out_0_8_1_port, P_OUT => lev_i_out_0_8_0_port)
                           ;
   PG_NETWORK_0_9 : PG_NET_56 port map( A => A(8), B => B(8), G_OUT => 
                           lev_i_out_0_9_1_port, P_OUT => lev_i_out_0_9_0_port)
                           ;
   PG_NETWORK_0_10 : PG_NET_55 port map( A => A(9), B => B(9), G_OUT => 
                           lev_i_out_0_10_1_port, P_OUT => 
                           lev_i_out_0_10_0_port);
   PG_NETWORK_0_11 : PG_NET_54 port map( A => A(10), B => B(10), G_OUT => 
                           lev_i_out_0_11_1_port, P_OUT => 
                           lev_i_out_0_11_0_port);
   PG_NETWORK_0_12 : PG_NET_53 port map( A => A(11), B => B(11), G_OUT => 
                           lev_i_out_0_12_1_port, P_OUT => 
                           lev_i_out_0_12_0_port);
   PG_NETWORK_0_13 : PG_NET_52 port map( A => A(12), B => B(12), G_OUT => 
                           lev_i_out_0_13_1_port, P_OUT => 
                           lev_i_out_0_13_0_port);
   PG_NETWORK_0_14 : PG_NET_51 port map( A => A(13), B => B(13), G_OUT => 
                           lev_i_out_0_14_1_port, P_OUT => 
                           lev_i_out_0_14_0_port);
   PG_NETWORK_0_15 : PG_NET_50 port map( A => A(14), B => B(14), G_OUT => 
                           lev_i_out_0_15_1_port, P_OUT => 
                           lev_i_out_0_15_0_port);
   PG_NETWORK_0_16 : PG_NET_49 port map( A => A(15), B => B(15), G_OUT => 
                           lev_i_out_0_16_1_port, P_OUT => 
                           lev_i_out_0_16_0_port);
   PG_NETWORK_0_17 : PG_NET_48 port map( A => A(16), B => B(16), G_OUT => 
                           lev_i_out_0_17_1_port, P_OUT => 
                           lev_i_out_0_17_0_port);
   PG_NETWORK_0_18 : PG_NET_47 port map( A => A(17), B => B(17), G_OUT => 
                           lev_i_out_0_18_1_port, P_OUT => 
                           lev_i_out_0_18_0_port);
   PG_NETWORK_0_19 : PG_NET_46 port map( A => A(18), B => B(18), G_OUT => 
                           lev_i_out_0_19_1_port, P_OUT => 
                           lev_i_out_0_19_0_port);
   PG_NETWORK_0_20 : PG_NET_45 port map( A => A(19), B => B(19), G_OUT => 
                           lev_i_out_0_20_1_port, P_OUT => 
                           lev_i_out_0_20_0_port);
   PG_NETWORK_0_21 : PG_NET_44 port map( A => A(20), B => B(20), G_OUT => 
                           lev_i_out_0_21_1_port, P_OUT => 
                           lev_i_out_0_21_0_port);
   PG_NETWORK_0_22 : PG_NET_43 port map( A => A(21), B => B(21), G_OUT => 
                           lev_i_out_0_22_1_port, P_OUT => 
                           lev_i_out_0_22_0_port);
   PG_NETWORK_0_23 : PG_NET_42 port map( A => A(22), B => B(22), G_OUT => 
                           lev_i_out_0_23_1_port, P_OUT => 
                           lev_i_out_0_23_0_port);
   PG_NETWORK_0_24 : PG_NET_41 port map( A => A(23), B => B(23), G_OUT => 
                           lev_i_out_0_24_1_port, P_OUT => 
                           lev_i_out_0_24_0_port);
   PG_NETWORK_0_25 : PG_NET_40 port map( A => A(24), B => B(24), G_OUT => 
                           lev_i_out_0_25_1_port, P_OUT => 
                           lev_i_out_0_25_0_port);
   PG_NETWORK_0_26 : PG_NET_39 port map( A => A(25), B => B(25), G_OUT => 
                           lev_i_out_0_26_1_port, P_OUT => 
                           lev_i_out_0_26_0_port);
   PG_NETWORK_0_27 : PG_NET_38 port map( A => A(26), B => B(26), G_OUT => 
                           lev_i_out_0_27_1_port, P_OUT => 
                           lev_i_out_0_27_0_port);
   PG_NETWORK_0_28 : PG_NET_37 port map( A => A(27), B => B(27), G_OUT => 
                           lev_i_out_0_28_1_port, P_OUT => 
                           lev_i_out_0_28_0_port);
   PG_NETWORK_0_29 : PG_NET_36 port map( A => A(28), B => B(28), G_OUT => 
                           lev_i_out_0_29_1_port, P_OUT => 
                           lev_i_out_0_29_0_port);
   PG_NETWORK_0_30 : PG_NET_35 port map( A => A(29), B => B(29), G_OUT => 
                           lev_i_out_0_30_1_port, P_OUT => 
                           lev_i_out_0_30_0_port);
   PG_NETWORK_0_31 : PG_NET_34 port map( A => A(30), B => B(30), G_OUT => 
                           lev_i_out_0_31_1_port, P_OUT => 
                           lev_i_out_0_31_0_port);
   PG_NETWORK_0_32 : PG_NET_33 port map( A => A(31), B => B(31), G_OUT => 
                           lev_i_out_0_32_1_port, P_OUT => 
                           lev_i_out_0_32_0_port);
   PG_NETWORK_0_33 : PG_NET_32 port map( A => A(32), B => B(32), G_OUT => 
                           lev_i_out_0_33_1_port, P_OUT => 
                           lev_i_out_0_33_0_port);
   PG_NETWORK_0_34 : PG_NET_31 port map( A => A(33), B => B(33), G_OUT => 
                           lev_i_out_0_34_1_port, P_OUT => 
                           lev_i_out_0_34_0_port);
   PG_NETWORK_0_35 : PG_NET_30 port map( A => A(34), B => B(34), G_OUT => 
                           lev_i_out_0_35_1_port, P_OUT => 
                           lev_i_out_0_35_0_port);
   PG_NETWORK_0_36 : PG_NET_29 port map( A => A(35), B => B(35), G_OUT => 
                           lev_i_out_0_36_1_port, P_OUT => 
                           lev_i_out_0_36_0_port);
   PG_NETWORK_0_37 : PG_NET_28 port map( A => A(36), B => B(36), G_OUT => 
                           lev_i_out_0_37_1_port, P_OUT => 
                           lev_i_out_0_37_0_port);
   PG_NETWORK_0_38 : PG_NET_27 port map( A => A(37), B => B(37), G_OUT => 
                           lev_i_out_0_38_1_port, P_OUT => 
                           lev_i_out_0_38_0_port);
   PG_NETWORK_0_39 : PG_NET_26 port map( A => A(38), B => B(38), G_OUT => 
                           lev_i_out_0_39_1_port, P_OUT => 
                           lev_i_out_0_39_0_port);
   PG_NETWORK_0_40 : PG_NET_25 port map( A => A(39), B => B(39), G_OUT => 
                           lev_i_out_0_40_1_port, P_OUT => 
                           lev_i_out_0_40_0_port);
   PG_NETWORK_0_41 : PG_NET_24 port map( A => A(40), B => B(40), G_OUT => 
                           lev_i_out_0_41_1_port, P_OUT => 
                           lev_i_out_0_41_0_port);
   PG_NETWORK_0_42 : PG_NET_23 port map( A => A(41), B => B(41), G_OUT => 
                           lev_i_out_0_42_1_port, P_OUT => 
                           lev_i_out_0_42_0_port);
   PG_NETWORK_0_43 : PG_NET_22 port map( A => A(42), B => B(42), G_OUT => 
                           lev_i_out_0_43_1_port, P_OUT => 
                           lev_i_out_0_43_0_port);
   PG_NETWORK_0_44 : PG_NET_21 port map( A => A(43), B => B(43), G_OUT => 
                           lev_i_out_0_44_1_port, P_OUT => 
                           lev_i_out_0_44_0_port);
   GNET1_1_2 : G_GENERAL_0 port map( PG_ik(1) => net102734, PG_ik(0) => 
                           lev_i_out_0_2_0_port, G_k_1j => lev_i_out_0_1_1_port
                           , G_ij => lev_i_out_1_2_1_port);
   PGNET1_1_4 : PG_GENERAL_0 port map( PG_ik(1) => lev_i_out_0_4_1_port, 
                           PG_ik(0) => lev_i_out_0_4_0_port, PG_k_1j(1) => 
                           lev_i_out_0_3_1_port, PG_k_1j(0) => 
                           lev_i_out_0_3_0_port, PG_ij(1) => 
                           lev_i_out_1_4_1_port, PG_ij(0) => 
                           lev_i_out_1_4_0_port);
   PGNET1_1_6 : PG_GENERAL_62 port map( PG_ik(1) => lev_i_out_0_6_1_port, 
                           PG_ik(0) => lev_i_out_0_6_0_port, PG_k_1j(1) => 
                           lev_i_out_0_5_1_port, PG_k_1j(0) => 
                           lev_i_out_0_5_0_port, PG_ij(1) => 
                           lev_i_out_1_6_1_port, PG_ij(0) => 
                           lev_i_out_1_6_0_port);
   PGNET1_1_8 : PG_GENERAL_61 port map( PG_ik(1) => lev_i_out_0_8_1_port, 
                           PG_ik(0) => lev_i_out_0_8_0_port, PG_k_1j(1) => 
                           lev_i_out_0_7_1_port, PG_k_1j(0) => 
                           lev_i_out_0_7_0_port, PG_ij(1) => 
                           lev_i_out_1_8_1_port, PG_ij(0) => 
                           lev_i_out_1_8_0_port);
   PGNET1_1_10 : PG_GENERAL_60 port map( PG_ik(1) => lev_i_out_0_10_1_port, 
                           PG_ik(0) => lev_i_out_0_10_0_port, PG_k_1j(1) => 
                           lev_i_out_0_9_1_port, PG_k_1j(0) => 
                           lev_i_out_0_9_0_port, PG_ij(1) => 
                           lev_i_out_1_10_1_port, PG_ij(0) => 
                           lev_i_out_1_10_0_port);
   PGNET1_1_12 : PG_GENERAL_59 port map( PG_ik(1) => lev_i_out_0_12_1_port, 
                           PG_ik(0) => lev_i_out_0_12_0_port, PG_k_1j(1) => 
                           lev_i_out_0_11_1_port, PG_k_1j(0) => 
                           lev_i_out_0_11_0_port, PG_ij(1) => 
                           lev_i_out_1_12_1_port, PG_ij(0) => 
                           lev_i_out_1_12_0_port);
   PGNET1_1_14 : PG_GENERAL_58 port map( PG_ik(1) => lev_i_out_0_14_1_port, 
                           PG_ik(0) => lev_i_out_0_14_0_port, PG_k_1j(1) => 
                           lev_i_out_0_13_1_port, PG_k_1j(0) => 
                           lev_i_out_0_13_0_port, PG_ij(1) => 
                           lev_i_out_1_14_1_port, PG_ij(0) => 
                           lev_i_out_1_14_0_port);
   PGNET1_1_16 : PG_GENERAL_57 port map( PG_ik(1) => lev_i_out_0_16_1_port, 
                           PG_ik(0) => lev_i_out_0_16_0_port, PG_k_1j(1) => 
                           lev_i_out_0_15_1_port, PG_k_1j(0) => 
                           lev_i_out_0_15_0_port, PG_ij(1) => 
                           lev_i_out_1_16_1_port, PG_ij(0) => 
                           lev_i_out_1_16_0_port);
   PGNET1_1_18 : PG_GENERAL_56 port map( PG_ik(1) => lev_i_out_0_18_1_port, 
                           PG_ik(0) => lev_i_out_0_18_0_port, PG_k_1j(1) => 
                           lev_i_out_0_17_1_port, PG_k_1j(0) => 
                           lev_i_out_0_17_0_port, PG_ij(1) => 
                           lev_i_out_1_18_1_port, PG_ij(0) => 
                           lev_i_out_1_18_0_port);
   PGNET1_1_20 : PG_GENERAL_55 port map( PG_ik(1) => lev_i_out_0_20_1_port, 
                           PG_ik(0) => lev_i_out_0_20_0_port, PG_k_1j(1) => 
                           lev_i_out_0_19_1_port, PG_k_1j(0) => 
                           lev_i_out_0_19_0_port, PG_ij(1) => 
                           lev_i_out_1_20_1_port, PG_ij(0) => 
                           lev_i_out_1_20_0_port, clk => clk);
   PGNET1_1_22 : PG_GENERAL_54 port map( PG_ik(1) => lev_i_out_0_22_1_port, 
                           PG_ik(0) => lev_i_out_0_22_0_port, PG_k_1j(1) => 
                           lev_i_out_0_21_1_port, PG_k_1j(0) => 
                           lev_i_out_0_21_0_port, PG_ij(1) => 
                           lev_i_out_1_22_1_port, PG_ij(0) => 
                           lev_i_out_1_22_0_port);
   PGNET1_1_24 : PG_GENERAL_53 port map( PG_ik(1) => lev_i_out_0_24_1_port, 
                           PG_ik(0) => lev_i_out_0_24_0_port, PG_k_1j(1) => 
                           lev_i_out_0_23_1_port, PG_k_1j(0) => 
                           lev_i_out_0_23_0_port, PG_ij(1) => 
                           lev_i_out_1_24_1_port, PG_ij(0) => 
                           lev_i_out_1_24_0_port);
   PGNET1_1_26 : PG_GENERAL_52 port map( PG_ik(1) => lev_i_out_0_26_1_port, 
                           PG_ik(0) => lev_i_out_0_26_0_port, PG_k_1j(1) => 
                           lev_i_out_0_25_1_port, PG_k_1j(0) => 
                           lev_i_out_0_25_0_port, PG_ij(1) => 
                           lev_i_out_1_26_1_port, PG_ij(0) => 
                           lev_i_out_1_26_0_port);
   PGNET1_1_28 : PG_GENERAL_51 port map( PG_ik(1) => lev_i_out_0_28_1_port, 
                           PG_ik(0) => lev_i_out_0_28_0_port, PG_k_1j(1) => 
                           lev_i_out_0_27_1_port, PG_k_1j(0) => 
                           lev_i_out_0_27_0_port, PG_ij(1) => 
                           lev_i_out_1_28_1_port, PG_ij(0) => 
                           lev_i_out_1_28_0_port);
   PGNET1_1_30 : PG_GENERAL_50 port map( PG_ik(1) => lev_i_out_0_30_1_port, 
                           PG_ik(0) => lev_i_out_0_30_0_port, PG_k_1j(1) => 
                           lev_i_out_0_29_1_port, PG_k_1j(0) => 
                           lev_i_out_0_29_0_port, PG_ij(1) => 
                           lev_i_out_1_30_1_port, PG_ij(0) => 
                           lev_i_out_1_30_0_port);
   PGNET1_1_32 : PG_GENERAL_49 port map( PG_ik(1) => lev_i_out_0_32_1_port, 
                           PG_ik(0) => lev_i_out_0_32_0_port, PG_k_1j(1) => 
                           lev_i_out_0_31_1_port, PG_k_1j(0) => 
                           lev_i_out_0_31_0_port, PG_ij(1) => 
                           lev_i_out_1_32_1_port, PG_ij(0) => 
                           lev_i_out_1_32_0_port);
   PGNET1_1_34 : PG_GENERAL_48 port map( PG_ik(1) => lev_i_out_0_34_1_port, 
                           PG_ik(0) => lev_i_out_0_34_0_port, PG_k_1j(1) => 
                           lev_i_out_0_33_1_port, PG_k_1j(0) => 
                           lev_i_out_0_33_0_port, PG_ij(1) => 
                           lev_i_out_1_34_1_port, PG_ij(0) => 
                           lev_i_out_1_34_0_port);
   PGNET1_1_36 : PG_GENERAL_47 port map( PG_ik(1) => lev_i_out_0_36_1_port, 
                           PG_ik(0) => lev_i_out_0_36_0_port, PG_k_1j(1) => 
                           lev_i_out_0_35_1_port, PG_k_1j(0) => 
                           lev_i_out_0_35_0_port, PG_ij(1) => 
                           lev_i_out_1_36_1_port, PG_ij(0) => 
                           lev_i_out_1_36_0_port);
   PGNET1_1_38 : PG_GENERAL_46 port map( PG_ik(1) => lev_i_out_0_38_1_port, 
                           PG_ik(0) => lev_i_out_0_38_0_port, PG_k_1j(1) => 
                           lev_i_out_0_37_1_port, PG_k_1j(0) => 
                           lev_i_out_0_37_0_port, PG_ij(1) => 
                           lev_i_out_1_38_1_port, PG_ij(0) => 
                           lev_i_out_1_38_0_port);
   PGNET1_1_40 : PG_GENERAL_45 port map( PG_ik(1) => lev_i_out_0_40_1_port, 
                           PG_ik(0) => lev_i_out_0_40_0_port, PG_k_1j(1) => 
                           lev_i_out_0_39_1_port, PG_k_1j(0) => 
                           lev_i_out_0_39_0_port, PG_ij(1) => 
                           lev_i_out_1_40_1_port, PG_ij(0) => 
                           lev_i_out_1_40_0_port);
   PGNET1_1_42 : PG_GENERAL_44 port map( PG_ik(1) => lev_i_out_0_42_1_port, 
                           PG_ik(0) => lev_i_out_0_42_0_port, PG_k_1j(1) => 
                           lev_i_out_0_41_1_port, PG_k_1j(0) => 
                           lev_i_out_0_41_0_port, PG_ij(1) => 
                           lev_i_out_1_42_1_port, PG_ij(0) => 
                           lev_i_out_1_42_0_port);
   PGNET1_1_44 : PG_GENERAL_43 port map( PG_ik(1) => lev_i_out_0_44_1_port, 
                           PG_ik(0) => lev_i_out_0_44_0_port, PG_k_1j(1) => 
                           lev_i_out_0_43_1_port, PG_k_1j(0) => 
                           lev_i_out_0_43_0_port, PG_ij(1) => 
                           lev_i_out_1_44_1_port, PG_ij(0) => 
                           lev_i_out_1_44_0_port);
   GNET_i_2_4_0 : G_GENERAL_16 port map( PG_ik(1) => lev_i_out_1_4_1_port, 
                           PG_ik(0) => lev_i_out_1_4_0_port, G_k_1j => 
                           lev_i_out_1_2_1_port, G_ij => n11, clk => clk);
   PGNET_i_2_8_0 : PG_GENERAL_32 port map( PG_ik(1) => lev_i_out_1_8_1_port, 
                           PG_ik(0) => lev_i_out_1_8_0_port, PG_k_1j(1) => 
                           lev_i_out_1_6_1_port, PG_k_1j(0) => 
                           lev_i_out_1_6_0_port, PG_ij(1) => 
                           lev_i_out_2_8_1_port, PG_ij(0) => 
                           lev_i_out_2_8_0_port);
   PGNET_i_2_12_0 : PG_GENERAL_31 port map( PG_ik(1) => lev_i_out_1_12_1_port, 
                           PG_ik(0) => lev_i_out_1_12_0_port, PG_k_1j(1) => 
                           lev_i_out_1_10_1_port, PG_k_1j(0) => 
                           lev_i_out_1_10_0_port, PG_ij(1) => 
                           lev_i_out_2_12_1_port, PG_ij(0) => 
                           lev_i_out_2_12_0_port);
   PGNET_i_2_16_0 : PG_GENERAL_30 port map( PG_ik(1) => lev_i_out_1_16_1_port, 
                           PG_ik(0) => lev_i_out_1_16_0_port, PG_k_1j(1) => 
                           lev_i_out_1_14_1_port, PG_k_1j(0) => 
                           lev_i_out_1_14_0_port, PG_ij(1) => 
                           lev_i_out_2_16_1_port, PG_ij(0) => 
                           lev_i_out_2_16_0_port, clk => clk);
   PGNET_i_2_20_0 : PG_GENERAL_29 port map( PG_ik(1) => lev_i_out_1_20_1_port, 
                           PG_ik(0) => lev_i_out_1_20_0_port, PG_k_1j(1) => 
                           lev_i_out_1_18_1_port, PG_k_1j(0) => 
                           lev_i_out_1_18_0_port, PG_ij(1) => 
                           lev_i_out_2_20_1_port, PG_ij(0) => 
                           lev_i_out_2_20_0_port, clk => clk);
   PGNET_i_2_24_0 : PG_GENERAL_28 port map( PG_ik(1) => lev_i_out_1_24_1_port, 
                           PG_ik(0) => lev_i_out_1_24_0_port, PG_k_1j(1) => 
                           lev_i_out_1_22_1_port, PG_k_1j(0) => 
                           lev_i_out_1_22_0_port, PG_ij(1) => 
                           lev_i_out_2_24_1_port, PG_ij(0) => 
                           lev_i_out_2_24_0_port);
   PGNET_i_2_28_0 : PG_GENERAL_27 port map( PG_ik(1) => lev_i_out_1_28_1_port, 
                           PG_ik(0) => lev_i_out_1_28_0_port, PG_k_1j(1) => 
                           lev_i_out_1_26_1_port, PG_k_1j(0) => 
                           lev_i_out_1_26_0_port, PG_ij(1) => n3, PG_ij(0) => 
                           lev_i_out_2_28_0_port);
   PGNET_i_2_32_0 : PG_GENERAL_26 port map( PG_ik(1) => lev_i_out_1_32_1_port, 
                           PG_ik(0) => lev_i_out_1_32_0_port, PG_k_1j(1) => 
                           lev_i_out_1_30_1_port, PG_k_1j(0) => 
                           lev_i_out_1_30_0_port, PG_ij(1) => 
                           lev_i_out_2_32_1_port, PG_ij(0) => 
                           lev_i_out_2_32_0_port);
   PGNET_i_2_36_0 : PG_GENERAL_25 port map( PG_ik(1) => lev_i_out_1_36_1_port, 
                           PG_ik(0) => lev_i_out_1_36_0_port, PG_k_1j(1) => 
                           lev_i_out_1_34_1_port, PG_k_1j(0) => 
                           lev_i_out_1_34_0_port, PG_ij(1) => 
                           lev_i_out_2_36_1_port, PG_ij(0) => 
                           lev_i_out_2_36_0_port);
   PGNET_i_2_40_0 : PG_GENERAL_24 port map( PG_ik(1) => lev_i_out_1_40_1_port, 
                           PG_ik(0) => lev_i_out_1_40_0_port, PG_k_1j(1) => 
                           lev_i_out_1_38_1_port, PG_k_1j(0) => 
                           lev_i_out_1_38_0_port, PG_ij(1) => 
                           lev_i_out_2_40_1_port, PG_ij(0) => 
                           lev_i_out_2_40_0_port);
   PGNET_i_2_44_0 : PG_GENERAL_23 port map( PG_ik(1) => lev_i_out_1_44_1_port, 
                           PG_ik(0) => lev_i_out_1_44_0_port, PG_k_1j(1) => 
                           lev_i_out_1_42_1_port, PG_k_1j(0) => 
                           lev_i_out_1_42_0_port, PG_ij(1) => 
                           lev_i_out_2_44_1_port, PG_ij(0) => 
                           lev_i_out_2_44_0_port);
   GNET_i_3_8_0 : G_GENERAL_15 port map( PG_ik(1) => lev_i_out_2_8_1_port, 
                           PG_ik(0) => lev_i_out_2_8_0_port, G_k_1j => n11, 
                           G_ij => n10);
   PGNET_i_3_16_0 : PG_GENERAL_17 port map( PG_ik(1) => lev_i_out_2_16_1_port, 
                           PG_ik(0) => lev_i_out_2_16_0_port, PG_k_1j(1) => 
                           lev_i_out_2_12_1_port, PG_k_1j(0) => 
                           lev_i_out_2_12_0_port, PG_ij(1) => 
                           lev_i_out_3_16_1_port, PG_ij(0) => 
                           lev_i_out_3_16_0_port, clk => clk);
   PGNET_i_3_24_0 : PG_GENERAL_16 port map( PG_ik(1) => lev_i_out_2_24_1_port, 
                           PG_ik(0) => lev_i_out_2_24_0_port, PG_k_1j(1) => 
                           lev_i_out_2_20_1_port, PG_k_1j(0) => 
                           lev_i_out_2_20_0_port, PG_ij(1) => 
                           lev_i_out_3_24_1_port, PG_ij(0) => 
                           lev_i_out_3_24_0_port);
   PGNET_i_3_32_0 : PG_GENERAL_15 port map( PG_ik(1) => lev_i_out_2_32_1_port, 
                           PG_ik(0) => lev_i_out_2_32_0_port, PG_k_1j(1) => n3,
                           PG_k_1j(0) => lev_i_out_2_28_0_port, PG_ij(1) => 
                           lev_i_out_3_32_1_port, PG_ij(0) => 
                           lev_i_out_3_32_0_port);
   PGNET_i_3_40_0 : PG_GENERAL_14 port map( PG_ik(1) => lev_i_out_2_40_1_port, 
                           PG_ik(0) => lev_i_out_2_40_0_port, PG_k_1j(1) => 
                           lev_i_out_2_36_1_port, PG_k_1j(0) => 
                           lev_i_out_2_36_0_port, PG_ij(1) => 
                           lev_i_out_3_40_1_port, PG_ij(0) => 
                           lev_i_out_3_40_0_port);
   GNET_i_4_16_0 : G_GENERAL_13 port map( PG_ik(1) => lev_i_out_3_16_1_port, 
                           PG_ik(0) => lev_i_out_3_16_0_port, G_k_1j => n10, 
                           G_ij => n9, clk => clk);
   PGNET_i_4_28_4 : PG_GENERAL_10 port map( PG_ik(1) => n3, PG_ik(0) => n15, 
                           PG_k_1j(1) => n14, PG_k_1j(0) => 
                           lev_i_out_3_24_0_port, PG_ij(1) => 
                           lev_i_out_4_28_1_port, PG_ij(0) => 
                           lev_i_out_4_28_0_port);
   PGNET_i_4_32_0 : PG_GENERAL_9 port map( PG_ik(1) => lev_i_out_3_32_1_port, 
                           PG_ik(0) => lev_i_out_3_32_0_port, PG_k_1j(1) => 
                           lev_i_out_3_24_1_port, PG_k_1j(0) => 
                           lev_i_out_3_24_0_port, PG_ij(1) => 
                           lev_i_out_4_32_1_port, PG_ij(0) => 
                           lev_i_out_4_32_0_port);
   PGNET_i_4_44_4 : PG_GENERAL_8 port map( PG_ik(1) => lev_i_out_2_44_1_port, 
                           PG_ik(0) => lev_i_out_2_44_0_port, PG_k_1j(1) => 
                           lev_i_out_3_40_1_port, PG_k_1j(0) => 
                           lev_i_out_3_40_0_port, PG_ij(1) => 
                           lev_i_out_4_44_1_port, PG_ij(0) => 
                           lev_i_out_4_44_0_port);
   GNET_i_5_20_12 : G_GENERAL_12 port map( PG_ik(1) => lev_i_out_2_20_1_port, 
                           PG_ik(0) => lev_i_out_2_20_0_port, G_k_1j => n9, 
                           G_ij => Co(5));
   GNET_i_5_24_8 : G_GENERAL_11 port map( PG_ik(1) => n14, PG_ik(0) => 
                           lev_i_out_3_24_0_port, G_k_1j => n9, G_ij => Co(6));
   GNET_i_5_28_4 : G_GENERAL_10 port map( PG_ik(1) => lev_i_out_4_28_1_port, 
                           PG_ik(0) => lev_i_out_4_28_0_port, G_k_1j => n9, 
                           G_ij => Co(7));
   GNET_i_5_32_0 : G_GENERAL_9 port map( PG_ik(1) => lev_i_out_4_32_1_port, 
                           PG_ik(0) => lev_i_out_4_32_0_port, G_k_1j => n9, 
                           G_ij => n8);
   GNET_i_6_36_28 : G_GENERAL_8 port map( PG_ik(1) => lev_i_out_2_36_1_port, 
                           PG_ik(0) => lev_i_out_2_36_0_port, G_k_1j => n8, 
                           G_ij => Co(9));
   GNET_i_6_40_24 : G_GENERAL_7 port map( PG_ik(1) => lev_i_out_3_40_1_port, 
                           PG_ik(0) => lev_i_out_3_40_0_port, G_k_1j => n8, 
                           G_ij => Co(10));
   GNET_i_6_44_20 : G_GENERAL_6 port map( PG_ik(1) => lev_i_out_4_44_1_port, 
                           PG_ik(0) => lev_i_out_4_44_0_port, G_k_1j => n8, 
                           G_ij => Co(11));
   U2 : CLKBUF_X1 port map( A => n8, Z => Co(8));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPround_SIG_width28_DW01_inc_1 is

   port( A : in std_logic_vector (24 downto 0);  SUM : out std_logic_vector (24
         downto 0));

end FPround_SIG_width28_DW01_inc_1;

architecture SYN_USE_DEFA_ARCH_NAME of FPround_SIG_width28_DW01_inc_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n6, n7, n11, n14, n16, n17, n18, n19, n23, n26, n28, n29, n31, 
      n35, n38, n40, n41, n50, n51, n52, n56, n57, n61, n62, n63, n68, n71, n73
      , n74, n76, n80, n83, n85, n86, n94, n95, n96, n97, n101, n105, n113, 
      n116, n123, n181, n182, n183, n184, n185, n186, n187, n188, n194, n196, 
      n197, n198, n200, n201, n203, n204, n207, n208, n209, n211, n212, n213, 
      n214, n218, n219, n220, n221, n222, n223, n224, n225, n226 : std_logic;

begin
   
   U154 : AND2_X1 port map( A1 => n28, A2 => n6, ZN => n181);
   U155 : XNOR2_X1 port map( A => n182, B => A(3), ZN => SUM(3));
   U156 : NAND2_X1 port map( A1 => n207, A2 => n200, ZN => n182);
   U157 : XOR2_X1 port map( A => n183, B => A(5), Z => SUM(5));
   U158 : NOR2_X1 port map( A1 => n212, A2 => n113, ZN => n183);
   U159 : XOR2_X1 port map( A => n184, B => A(6), Z => SUM(6));
   U160 : NOR2_X1 port map( A1 => n212, A2 => n197, ZN => n184);
   U161 : XOR2_X1 port map( A => n185, B => A(7), Z => SUM(7));
   U162 : NOR2_X1 port map( A1 => n212, A2 => n101, ZN => n185);
   U163 : XNOR2_X1 port map( A => n186, B => A(9), ZN => SUM(9));
   U164 : NAND2_X1 port map( A1 => n94, A2 => A(8), ZN => n186);
   U165 : XNOR2_X1 port map( A => n187, B => A(11), ZN => SUM(11));
   U166 : NAND2_X1 port map( A1 => n94, A2 => n80, ZN => n187);
   U167 : XNOR2_X1 port map( A => n188, B => A(13), ZN => SUM(13));
   U168 : NAND2_X1 port map( A1 => n68, A2 => n94, ZN => n188);
   U179 : XNOR2_X1 port map( A => n194, B => A(23), ZN => SUM(23));
   U180 : NAND2_X1 port map( A1 => n214, A2 => n11, ZN => n194);
   U183 : INV_X1 port map( A => n211, ZN => n74);
   U185 : NOR2_X1 port map( A1 => n19, A2 => n7, ZN => n6);
   U186 : NOR2_X1 port map( A1 => n201, A2 => n38, ZN => n35);
   U187 : NOR2_X1 port map( A1 => n86, A2 => n83, ZN => n80);
   U188 : NOR2_X1 port map( A1 => n29, A2 => n26, ZN => n23);
   U189 : INV_X1 port map( A => n28, ZN => n29);
   U191 : NOR2_X1 port map( A1 => n74, A2 => n62, ZN => n61);
   U192 : NOR2_X1 port map( A1 => n74, A2 => n71, ZN => n68);
   U193 : NOR2_X1 port map( A1 => n17, A2 => n14, ZN => n11);
   U194 : NAND2_X1 port map( A1 => n28, A2 => n18, ZN => n17);
   U195 : INV_X1 port map( A => n19, ZN => n18);
   U197 : NAND2_X1 port map( A1 => n73, A2 => n51, ZN => n50);
   U198 : NOR2_X1 port map( A1 => n62, A2 => n52, ZN => n51);
   U199 : NAND2_X1 port map( A1 => A(14), A2 => A(15), ZN => n52);
   U201 : NAND2_X1 port map( A1 => A(18), A2 => A(19), ZN => n31);
   U203 : NAND2_X1 port map( A1 => A(10), A2 => A(11), ZN => n76);
   U205 : NAND2_X1 port map( A1 => A(2), A2 => A(3), ZN => n116);
   U206 : XOR2_X1 port map( A => n213, B => A(16), Z => SUM(16));
   U207 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n41);
   U211 : INV_X1 port map( A => n86, ZN => n85);
   U216 : INV_X1 port map( A => n201, ZN => n40);
   U221 : INV_X1 port map( A => n17, ZN => n16);
   U222 : INV_X1 port map( A => A(18), ZN => n38);
   U223 : INV_X1 port map( A => A(20), ZN => n26);
   U224 : INV_X1 port map( A => A(10), ZN => n83);
   U225 : INV_X1 port map( A => A(22), ZN => n14);
   U226 : INV_X1 port map( A => A(12), ZN => n71);
   U227 : INV_X1 port map( A => A(4), ZN => n113);
   U228 : XOR2_X1 port map( A => n212, B => n113, Z => SUM(4));
   U229 : NAND2_X1 port map( A1 => A(4), A2 => A(5), ZN => n105);
   U231 : XOR2_X1 port map( A => n94, B => A(8), Z => SUM(8));
   U232 : NOR2_X1 port map( A1 => n74, A2 => n57, ZN => n56);
   U233 : NAND2_X1 port map( A1 => n63, A2 => A(14), ZN => n57);
   U234 : INV_X1 port map( A => n62, ZN => n63);
   U235 : NAND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n123);
   U236 : NAND2_X1 port map( A1 => A(20), A2 => A(21), ZN => n19);
   U237 : NAND2_X1 port map( A1 => n223, A2 => A(6), ZN => n101);
   U239 : NAND2_X1 port map( A1 => A(22), A2 => A(23), ZN => n7);
   U240 : NAND2_X1 port map( A1 => n204, A2 => n208, ZN => n95);
   U241 : NOR2_X1 port map( A1 => n105, A2 => n97, ZN => n96);
   U242 : NAND2_X1 port map( A1 => A(6), A2 => A(7), ZN => n97);
   U243 : XOR2_X1 port map( A => n207, B => n200, Z => SUM(2));
   U244 : INV_X1 port map( A => n224, ZN => SUM(0));
   U245 : XOR2_X1 port map( A => A(1), B => n224, Z => SUM(1));
   U184 : AND2_X1 port map( A1 => n1, A2 => n181, ZN => SUM(24));
   U169 : XOR2_X1 port map( A => n196, B => A(14), Z => SUM(14));
   U170 : AND2_X1 port map( A1 => n94, A2 => n61, ZN => n196);
   U177 : INV_X1 port map( A => n223, ZN => n197);
   U178 : XOR2_X1 port map( A => n198, B => A(21), Z => SUM(21));
   U181 : AND2_X1 port map( A1 => n213, A2 => n23, ZN => n198);
   U190 : CLKBUF_X1 port map( A => A(2), Z => n200);
   U200 : NAND2_X1 port map( A1 => A(16), A2 => A(17), ZN => n201);
   U220 : XNOR2_X1 port map( A => n203, B => n14, ZN => SUM(22));
   U246 : AND2_X1 port map( A1 => n214, A2 => n16, ZN => n203);
   U248 : NOR2_X1 port map( A1 => n105, A2 => n97, ZN => n204);
   U250 : AND2_X1 port map( A1 => A(1), A2 => n224, ZN => n207);
   U251 : NOR2_X1 port map( A1 => n116, A2 => n123, ZN => n208);
   U252 : NOR2_X2 port map( A1 => n209, A2 => n50, ZN => n213);
   U253 : NAND2_X1 port map( A1 => n96, A2 => n208, ZN => n209);
   U255 : NOR2_X1 port map( A1 => n86, A2 => n76, ZN => n211);
   U256 : NOR2_X1 port map( A1 => n86, A2 => n76, ZN => n73);
   U257 : OR2_X1 port map( A1 => n116, A2 => n123, ZN => n212);
   U258 : NOR2_X1 port map( A1 => n50, A2 => n209, ZN => n214);
   U259 : NOR2_X1 port map( A1 => n50, A2 => n95, ZN => n1);
   U247 : NOR2_X1 port map( A1 => n41, A2 => n31, ZN => n28);
   U208 : NAND2_X1 port map( A1 => A(8), A2 => A(9), ZN => n86);
   U230 : NAND2_X1 port map( A1 => A(12), A2 => A(13), ZN => n62);
   U171 : BUF_X1 port map( A => A(0), Z => n224);
   U172 : XOR2_X1 port map( A => n218, B => A(15), Z => SUM(15));
   U173 : AND2_X1 port map( A1 => n94, A2 => n56, ZN => n218);
   U174 : XOR2_X1 port map( A => n219, B => A(19), Z => SUM(19));
   U175 : AND2_X1 port map( A1 => n213, A2 => n35, ZN => n219);
   U176 : INV_X1 port map( A => n209, ZN => n94);
   U182 : XNOR2_X1 port map( A => n220, B => n71, ZN => SUM(12));
   U196 : AND2_X1 port map( A1 => n94, A2 => n211, ZN => n220);
   U202 : XOR2_X1 port map( A => n221, B => A(17), Z => SUM(17));
   U204 : AND2_X1 port map( A1 => n213, A2 => A(16), ZN => n221);
   U209 : XNOR2_X1 port map( A => n222, B => n83, ZN => SUM(10));
   U210 : AND2_X1 port map( A1 => n94, A2 => n85, ZN => n222);
   U212 : AND2_X1 port map( A1 => A(4), A2 => A(5), ZN => n223);
   U213 : XNOR2_X1 port map( A => n225, B => n26, ZN => SUM(20));
   U214 : AND2_X1 port map( A1 => n213, A2 => n28, ZN => n225);
   U215 : XNOR2_X1 port map( A => n226, B => n38, ZN => SUM(18));
   U217 : AND2_X1 port map( A1 => n213, A2 => n40, ZN => n226);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (63 downto 0);  Cout : out std_logic;  clk : in 
         std_logic);

end P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRS_X2
      port( D, CK, RN, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic_vector
            (15 downto 0);  S : out std_logic_vector (63 downto 0);  clk : in 
            std_logic);
   end component;
   
   component CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (16 downto 0);  clk : in std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n151, n152, carry_out_11_port, carry_out_10_port, carry_out_9_port, 
      carry_out_8_port, carry_out_7_port, carry_out_6_port, carry_out_5_port, 
      n6, n14, n24, n25, n26, n29, n32, n36, n2, n3, n4, n5, n8, n20, n22, n30,
      n37, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52
      , n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n154, n155, n156, n157, n158, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n217, n220, n221, n_1448, n_1449, n_1450, n_1451, 
      n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, 
      n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, 
      n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, 
      n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, 
      n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, 
      n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, 
      n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, 
      n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523 : 
      std_logic;

begin
   
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';
   n8 <= '0';
   n20 <= '0';
   n22 <= '0';
   n30 <= '0';
   n37 <= '0';
   n39 <= '0';
   n40 <= '0';
   n41 <= '0';
   n42 <= '0';
   n43 <= '0';
   n44 <= '0';
   n45 <= '0';
   n46 <= '0';
   n47 <= '0';
   n48 <= '0';
   n49 <= '0';
   n50 <= '0';
   n51 <= '0';
   n52 <= '0';
   n53 <= '0';
   n54 <= '0';
   n55 <= '0';
   n56 <= '0';
   n57 <= '0';
   n58 <= '0';
   n59 <= '0';
   n60 <= '0';
   n61 <= '0';
   n62 <= '0';
   n63 <= '0';
   n64 <= '0';
   n65 <= '0';
   n66 <= '0';
   n67 <= '0';
   n68 <= '0';
   n69 <= '0';
   n70 <= '0';
   n71 <= '0';
   n72 <= '0';
   n73 <= '0';
   n74 <= '0';
   n75 <= '0';
   n76 <= '0';
   n77 <= '0';
   n78 <= '0';
   n79 <= '0';
   n80 <= '0';
   n81 <= '0';
   n82 <= '0';
   n83 <= '0';
   n84 <= '0';
   n85 <= '0';
   n86 <= '0';
   n87 <= '0';
   n88 <= '0';
   n89 <= '0';
   n90 <= '0';
   n91 <= '0';
   n92 <= '0';
   n93 <= '0';
   n94 <= '0';
   n95 <= '0';
   n96 <= '0';
   n97 <= '0';
   n98 <= '0';
   n99 <= '0';
   n100 <= '0';
   n101 <= '0';
   n102 <= '0';
   n103 <= '0';
   n104 <= '0';
   n105 <= '0';
   n106 <= '0';
   n107 <= '0';
   n108 <= '0';
   n109 <= '0';
   n110 <= '0';
   n111 <= '0';
   n112 <= '0';
   n113 <= '0';
   n114 <= '0';
   n115 <= '0';
   n116 <= '0';
   n117 <= '0';
   n118 <= '0';
   n119 <= '0';
   n120 <= '0';
   n121 <= '0';
   n122 <= '0';
   n123 <= '0';
   n124 <= '0';
   n125 <= '0';
   n126 <= '0';
   n127 <= '0';
   n128 <= '0';
   n129 <= '0';
   n130 <= '0';
   n131 <= '0';
   n132 <= '0';
   n133 <= '0';
   n134 <= '0';
   n135 <= '0';
   n136 <= '0';
   n137 <= '0';
   n138 <= '0';
   n139 <= '0';
   n140 <= '0';
   n141 <= '0';
   n142 <= '0';
   n143 <= '0';
   n144 <= '0';
   n145 <= '0';
   n146 <= '0';
   n147 <= '0';
   n148 <= '0';
   n149 <= '0';
   n150 <= '0';
   U10 : CLKBUF_X1 port map( A => n192, Z => n14);
   U11 : CLKBUF_X1 port map( A => n196, Z => n24);
   n152 <= '0';
   n151 <= '0';
   U17 : CLKBUF_X1 port map( A => n190, Z => n154);
   U19 : CLKBUF_X1 port map( A => n204, Z => n158);
   MY_CLK_r_REG353_S2 : DFF_X1 port map( D => A(43), CK => clk, Q => n214, QN 
                           => n_1448);
   MY_CLK_r_REG298_S2 : DFF_X1 port map( D => A(33), CK => clk, Q => n213, QN 
                           => n_1449);
   MY_CLK_r_REG282_S2 : DFF_X1 port map( D => A(30), CK => clk, Q => n211, QN 
                           => n_1450);
   MY_CLK_r_REG273_S2 : DFF_X1 port map( D => A(28), CK => clk, Q => n209, QN 
                           => n_1451);
   MY_CLK_r_REG257_S2 : DFF_X1 port map( D => A(27), CK => clk, Q => n208, QN 
                           => n_1452);
   MY_CLK_r_REG260_S2 : DFF_X1 port map( D => A(26), CK => clk, Q => n207, QN 
                           => n_1453);
   MY_CLK_r_REG263_S2 : DFF_X1 port map( D => A(25), CK => clk, Q => n206, QN 
                           => n_1454);
   MY_CLK_r_REG266_S2 : DFF_X1 port map( D => A(24), CK => clk, Q => n205, QN 
                           => n_1455);
   MY_CLK_r_REG414_S2 : DFF_X1 port map( D => A(22), CK => clk, Q => n203, QN 
                           => n_1456);
   MY_CLK_r_REG434_S2 : DFF_X1 port map( D => A(21), CK => clk, Q => n202, QN 
                           => n_1457);
   MY_CLK_r_REG444_S2 : DFF_X1 port map( D => A(20), CK => clk, Q => n201, QN 
                           => n_1458);
   MY_CLK_r_REG297_S2 : DFF_X1 port map( D => B(34), CK => clk, Q => n200, QN 
                           => n_1459);
   MY_CLK_r_REG293_S2 : DFF_X1 port map( D => B(33), CK => clk, Q => n199, QN 
                           => n_1460);
   MY_CLK_r_REG281_S2 : DFF_X1 port map( D => B(31), CK => clk, Q => n198, QN 
                           => n_1461);
   MY_CLK_r_REG278_S2 : DFF_X1 port map( D => B(30), CK => clk, Q => n197, QN 
                           => n_1462);
   MY_CLK_r_REG274_S2 : DFF_X1 port map( D => B(29), CK => clk, Q => n196, QN 
                           => n_1463);
   MY_CLK_r_REG201_S2 : DFF_X1 port map( D => B(28), CK => clk, Q => n195, QN 
                           => n_1464);
   MY_CLK_r_REG259_S2 : DFF_X1 port map( D => B(27), CK => clk, Q => n194, QN 
                           => n_1465);
   MY_CLK_r_REG262_S2 : DFF_X1 port map( D => B(26), CK => clk, Q => n193, QN 
                           => n_1466);
   MY_CLK_r_REG265_S2 : DFF_X1 port map( D => B(25), CK => clk, Q => n192, QN 
                           => n_1467);
   MY_CLK_r_REG269_S2 : DFF_X1 port map( D => B(24), CK => clk, Q => n191, QN 
                           => n_1468);
   MY_CLK_r_REG413_S2 : DFF_X1 port map( D => B(23), CK => clk, Q => n190, QN 
                           => n_1469);
   MY_CLK_r_REG435_S2 : DFF_X1 port map( D => B(22), CK => clk, Q => n189, QN 
                           => n_1470);
   MY_CLK_r_REG443_S2 : DFF_X1 port map( D => B(21), CK => clk, Q => n188, QN 
                           => n_1471);
   MY_CLK_r_REG459_S2 : DFF_X1 port map( D => B(20), CK => clk, Q => n187, QN 
                           => n_1472);
   MY_CLK_r_REG283_S2 : DFF_X1 port map( D => A(31), CK => clk, Q => n212, QN 
                           => n_1473);
   MY_CLK_r_REG270_S2 : DFF_X1 port map( D => A(23), CK => clk, Q => n204, QN 
                           => n_1474);
   U13 : CLKBUF_X1 port map( A => n197, Z => n32);
   U7 : CLKBUF_X1 port map( A => n189, Z => n6);
   U30 : CLKBUF_X1 port map( A => n193, Z => n29);
   U27 : CLKBUF_X1 port map( A => A(35), Z => n26);
   U29 : BUF_X1 port map( A => A(36), Z => n156);
   U8 : BUF_X1 port map( A => n188, Z => n217);
   U12 : BUF_X1 port map( A => n202, Z => n36);
   U14 : CLKBUF_X1 port map( A => n198, Z => n25);
   U18 : CLKBUF_X1 port map( A => A(37), Z => n155);
   U20 : CLKBUF_X1 port map( A => A(39), Z => n157);
   CARRY_GEN_INST : CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4 port map( A(63) => 
                           n2, A(62) => n3, A(61) => n4, A(60) => n5, A(59) => 
                           n8, A(58) => n20, A(57) => n22, A(56) => n30, A(55) 
                           => n37, A(54) => n39, A(53) => n40, A(52) => n41, 
                           A(51) => n42, A(50) => n43, A(49) => n44, A(48) => 
                           n45, A(47) => n46, A(46) => n47, A(45) => n48, A(44)
                           => n49, A(43) => n214, A(42) => A(42), A(41) => 
                           A(41), A(40) => A(40), A(39) => A(39), A(38) => 
                           A(38), A(37) => A(37), A(36) => A(36), A(35) => 
                           A(35), A(34) => A(34), A(33) => n213, A(32) => A(32)
                           , A(31) => n212, A(30) => n211, A(29) => n210, A(28)
                           => n209, A(27) => n208, A(26) => n207, A(25) => n206
                           , A(24) => n205, A(23) => n204, A(22) => n203, A(21)
                           => n202, A(20) => n201, A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(63) => n50, B(62) => n51, 
                           B(61) => n52, B(60) => n53, B(59) => n54, B(58) => 
                           n55, B(57) => n56, B(56) => n57, B(55) => n58, B(54)
                           => n59, B(53) => n60, B(52) => n61, B(51) => n62, 
                           B(50) => n63, B(49) => n64, B(48) => n65, B(47) => 
                           n66, B(46) => n67, B(45) => n68, B(44) => n69, B(43)
                           => B(43), B(42) => B(42), B(41) => B(41), B(40) => 
                           B(40), B(39) => B(39), B(38) => B(38), B(37) => 
                           B(37), B(36) => B(36), B(35) => B(35), B(34) => n200
                           , B(33) => n199, B(32) => B(32), B(31) => n198, 
                           B(30) => n197, B(29) => n196, B(28) => n195, B(27) 
                           => n194, B(26) => n193, B(25) => n192, B(24) => n191
                           , B(23) => n190, B(22) => n189, B(21) => n188, B(20)
                           => n187, B(19) => B(19), B(18) => B(18), B(17) => 
                           B(17), B(16) => B(16), B(15) => B(15), B(14) => 
                           B(14), B(13) => B(13), B(12) => B(12), B(11) => 
                           B(11), B(10) => B(10), B(9) => B(9), B(8) => B(8), 
                           B(7) => B(7), B(6) => B(6), B(5) => B(5), B(4) => 
                           B(4), B(3) => B(3), B(2) => B(2), B(1) => n151, B(0)
                           => B(0), Cin => n152, Co(16) => n_1475, Co(15) => 
                           n_1476, Co(14) => n_1477, Co(13) => n_1478, Co(12) 
                           => n_1479, Co(11) => carry_out_11_port, Co(10) => 
                           carry_out_10_port, Co(9) => carry_out_9_port, Co(8) 
                           => carry_out_8_port, Co(7) => carry_out_7_port, 
                           Co(6) => carry_out_6_port, Co(5) => carry_out_5_port
                           , Co(4) => n_1480, Co(3) => n_1481, Co(2) => n_1482,
                           Co(1) => n_1483, Co(0) => n_1484, clk => clk);
   SUM_GEN_INST : SUM_GENERATOR_NBIT_PER_BLOCK4_NBLOCKS16 port map( A(63) => 
                           n70, A(62) => n71, A(61) => n72, A(60) => n73, A(59)
                           => n74, A(58) => n75, A(57) => n76, A(56) => n77, 
                           A(55) => n78, A(54) => n79, A(53) => n80, A(52) => 
                           n81, A(51) => n82, A(50) => n83, A(49) => n84, A(48)
                           => n85, A(47) => A(47), A(46) => A(46), A(45) => 
                           A(45), A(44) => A(44), A(43) => n214, A(42) => A(42)
                           , A(41) => A(41), A(40) => A(40), A(39) => n157, 
                           A(38) => A(38), A(37) => n155, A(36) => n156, A(35) 
                           => n26, A(34) => A(34), A(33) => n213, A(32) => 
                           A(32), A(31) => n212, A(30) => n211, A(29) => n210, 
                           A(28) => n209, A(27) => n208, A(26) => n207, A(25) 
                           => n206, A(24) => n205, A(23) => n158, A(22) => n203
                           , A(21) => n36, A(20) => n201, A(19) => n86, A(18) 
                           => n87, A(17) => n88, A(16) => n89, A(15) => n90, 
                           A(14) => n91, A(13) => n92, A(12) => n93, A(11) => 
                           n94, A(10) => n95, A(9) => n96, A(8) => n97, A(7) =>
                           n98, A(6) => n99, A(5) => n100, A(4) => n101, A(3) 
                           => n102, A(2) => n103, A(1) => n104, A(0) => n105, 
                           B(63) => n106, B(62) => n107, B(61) => n108, B(60) 
                           => n109, B(59) => n110, B(58) => n111, B(57) => n112
                           , B(56) => n113, B(55) => n114, B(54) => n115, B(53)
                           => n116, B(52) => n117, B(51) => n118, B(50) => n119
                           , B(49) => n120, B(48) => n121, B(47) => B(47), 
                           B(46) => B(46), B(45) => B(45), B(44) => B(44), 
                           B(43) => B(43), B(42) => B(42), B(41) => B(41), 
                           B(40) => B(40), B(39) => B(39), B(38) => B(38), 
                           B(37) => B(37), B(36) => B(36), B(35) => B(35), 
                           B(34) => n200, B(33) => n199, B(32) => B(32), B(31) 
                           => n25, B(30) => n32, B(29) => n24, B(28) => n195, 
                           B(27) => n220, B(26) => n29, B(25) => n14, B(24) => 
                           n191, B(23) => n154, B(22) => n6, B(21) => n217, 
                           B(20) => n187, B(19) => n122, B(18) => n123, B(17) 
                           => n124, B(16) => n125, B(15) => n126, B(14) => n127
                           , B(13) => n128, B(12) => n129, B(11) => n130, B(10)
                           => n131, B(9) => n132, B(8) => n133, B(7) => n134, 
                           B(6) => n135, B(5) => n136, B(4) => n137, B(3) => 
                           n138, B(2) => n139, B(1) => n140, B(0) => n141, 
                           Ci(15) => n142, Ci(14) => n143, Ci(13) => n144, 
                           Ci(12) => n145, Ci(11) => carry_out_11_port, Ci(10) 
                           => carry_out_10_port, Ci(9) => carry_out_9_port, 
                           Ci(8) => carry_out_8_port, Ci(7) => carry_out_7_port
                           , Ci(6) => carry_out_6_port, Ci(5) => 
                           carry_out_5_port, Ci(4) => n146, Ci(3) => n147, 
                           Ci(2) => n148, Ci(1) => n149, Ci(0) => n150, S(63) 
                           => n_1485, S(62) => n_1486, S(61) => n_1487, S(60) 
                           => n_1488, S(59) => n_1489, S(58) => n_1490, S(57) 
                           => n_1491, S(56) => n_1492, S(55) => n_1493, S(54) 
                           => n_1494, S(53) => n_1495, S(52) => n_1496, S(51) 
                           => n_1497, S(50) => n_1498, S(49) => n_1499, S(48) 
                           => n_1500, S(47) => S(47), S(46) => S(46), S(45) => 
                           S(45), S(44) => S(44), S(43) => S(43), S(42) => 
                           S(42), S(41) => S(41), S(40) => S(40), S(39) => 
                           S(39), S(38) => S(38), S(37) => S(37), S(36) => 
                           S(36), S(35) => S(35), S(34) => S(34), S(33) => 
                           S(33), S(32) => S(32), S(31) => S(31), S(30) => 
                           S(30), S(29) => S(29), S(28) => S(28), S(27) => 
                           S(27), S(26) => S(26), S(25) => S(25), S(24) => 
                           S(24), S(23) => S(23), S(22) => S(22), S(21) => 
                           n_1501, S(20) => n_1502, S(19) => n_1503, S(18) => 
                           n_1504, S(17) => n_1505, S(16) => n_1506, S(15) => 
                           n_1507, S(14) => n_1508, S(13) => n_1509, S(12) => 
                           n_1510, S(11) => n_1511, S(10) => n_1512, S(9) => 
                           n_1513, S(8) => n_1514, S(7) => n_1515, S(6) => 
                           n_1516, S(5) => n_1517, S(4) => n_1518, S(3) => 
                           n_1519, S(2) => n_1520, S(1) => n_1521, S(0) => 
                           n_1522, clk => clk);
   MY_CLK_r_REG277_S2 : DFFRS_X2 port map( D => A(29), CK => clk, RN => n221, 
                           SN => n221, Q => n210, QN => n_1523);
   U6 : CLKBUF_X1 port map( A => n194, Z => n220);
   n221 <= '1';

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U1 : XNOR2_X1 port map( A => B, B => n2, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XNOR2_X1 port map( A => n1, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U5 : INV_X1 port map( A => B, ZN => n1);
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U4 : INV_X1 port map( A => B, ZN => n4);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n8, n9 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n9, A2 => n8, ZN => Co);
   U2 : XOR2_X1 port map( A => n6, B => n5, Z => S);
   MY_CLK_r_REG354_S2 : DFF_X1 port map( D => A, CK => clk, Q => n6, QN => n9);
   MY_CLK_r_REG338_S2 : DFF_X1 port map( D => B, CK => clk, Q => n5, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n8, n_1532 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => n6, ZN => S);
   U4 : INV_X1 port map( A => B, ZN => n4);
   U2 : NOR2_X1 port map( A1 => n8, A2 => n6, ZN => Co);
   MY_CLK_r_REG339_S2 : DFF_X1 port map( D => n4, CK => clk, Q => n6, QN => 
                           n_1532);
   MY_CLK_r_REG337_S2 : DFF_X1 port map( D => A, CK => clk, Q => n5, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5, n7, n_1534 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => n7, ZN => S);
   MY_CLK_r_REG332_S2 : DFF_X1 port map( D => B, CK => clk, Q => n3, QN => n7);
   MY_CLK_r_REG340_S2 : DFF_X1 port map( D => A, CK => clk, Q => n5, QN => 
                           n_1534);
   U2 : AND2_X1 port map( A1 => n5, A2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n3, n4, n8, n_1536 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n3, B => n4, ZN => S);
   U1 : NOR2_X1 port map( A1 => n8, A2 => n4, ZN => Co);
   U2 : INV_X1 port map( A => B, ZN => n6);
   MY_CLK_r_REG329_S2 : DFF_X1 port map( D => n6, CK => clk, Q => n4, QN => 
                           n_1536);
   MY_CLK_r_REG333_S2 : DFF_X1 port map( D => A, CK => clk, Q => n3, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5, n7, n_1538 : std_logic;

begin
   
   U2 : AND2_X1 port map( A1 => n3, A2 => n5, ZN => Co);
   MY_CLK_r_REG328_S2 : DFF_X1 port map( D => A, CK => clk, Q => n5, QN => 
                           n_1538);
   MY_CLK_r_REG319_S2 : DFF_X1 port map( D => B, CK => clk, Q => n3, QN => n7);
   U1 : XNOR2_X1 port map( A => n5, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5, n7, n8, n_1540 : std_logic;

begin
   
   U1 : INV_X1 port map( A => B, ZN => n3);
   U2 : NOR2_X2 port map( A1 => n7, A2 => n5, ZN => Co);
   MY_CLK_r_REG321_S2 : DFF_X1 port map( D => n3, CK => clk, Q => n5, QN => n8)
                           ;
   MY_CLK_r_REG320_S2 : DFF_X1 port map( D => A, CK => clk, Q => n_1540, QN => 
                           n7);
   U3 : XNOR2_X1 port map( A => n7, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5, n7, n_1542 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => n7, ZN => S);
   MY_CLK_r_REG322_S2 : DFF_X1 port map( D => A, CK => clk, Q => n5, QN => 
                           n_1542);
   MY_CLK_r_REG308_S2 : DFF_X1 port map( D => B, CK => clk, Q => n3, QN => n7);
   U1 : AND2_X2 port map( A1 => n5, A2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n4, n8, n9, n_1544 : std_logic;

begin
   
   U2 : INV_X1 port map( A => B, ZN => n6);
   U1 : NOR2_X2 port map( A1 => n8, A2 => n4, ZN => Co);
   MY_CLK_r_REG310_S2 : DFF_X1 port map( D => n6, CK => clk, Q => n4, QN => n9)
                           ;
   MY_CLK_r_REG309_S2 : DFF_X1 port map( D => A, CK => clk, Q => n_1544, QN => 
                           n8);
   U3 : XNOR2_X1 port map( A => n8, B => n9, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n3, n5, n7, n_1546 : std_logic;

begin
   
   MY_CLK_r_REG311_S2 : DFF_X1 port map( D => A, CK => clk, Q => n5, QN => n7);
   MY_CLK_r_REG302_S2 : DFF_X1 port map( D => B, CK => clk, Q => n3, QN => 
                           n_1546);
   U1 : XNOR2_X1 port map( A => n7, B => n3, ZN => S);
   U2 : AND2_X2 port map( A1 => n5, A2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => Co);
   U1 : XOR2_X1 port map( A => A, B => B, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n_1548, n_1549 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n3);
   MY_CLK_r_REG299_S2 : DFF_X1 port map( D => A, CK => clk, Q => n7, QN => 
                           n_1548);
   MY_CLK_r_REG292_S2 : DFF_X1 port map( D => n3, CK => clk, Q => n6, QN => 
                           n_1549);
   U5 : OAI21_X1 port map( B1 => Ci, B2 => B, A => A, ZN => n5);
   U4 : XNOR2_X2 port map( A => n7, B => n6, ZN => S);
   U2 : NAND2_X1 port map( A1 => B, A2 => Ci, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27308, net27309, net27310, net34232, n1, n5, n6, n7, n_1550, 
      n_1551, n_1552 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : INV_X1 port map( A => B, ZN => net27309);
   U4 : CLKBUF_X1 port map( A => A, Z => net34232);
   U5 : OAI21_X1 port map( B1 => net34232, B2 => B, A => Ci, ZN => net27310);
   U6 : INV_X1 port map( A => net34232, ZN => net27308);
   MY_CLK_r_REG284_S2 : DFF_X1 port map( D => net27309, CK => clk, Q => n7, QN 
                           => n_1550);
   MY_CLK_r_REG291_S2 : DFF_X1 port map( D => net27308, CK => clk, Q => n6, QN 
                           => n_1551);
   MY_CLK_r_REG285_S2 : DFF_X1 port map( D => net27310, CK => clk, Q => n5, QN 
                           => n_1552);
   U8 : OAI21_X2 port map( B1 => n6, B2 => n7, A => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27312, net27313, n2 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net27312);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net27313);
   U7 : NAND2_X1 port map( A1 => net27313, A2 => net27312, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27315, net27316, net27317, net31457, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U4 : OAI21_X1 port map( B1 => net31457, B2 => B, A => Ci, ZN => net27317);
   U5 : INV_X1 port map( A => B, ZN => net27316);
   U6 : OAI21_X1 port map( B1 => net27315, B2 => net27316, A => net27317, ZN =>
                           Co);
   U7 : INV_X1 port map( A => net31457, ZN => net27315);
   U3 : CLKBUF_X1 port map( A => A, Z => net31457);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n2, B => A, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => Ci, ZN => n2);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U1 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27323, net27324, net27325, n2 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => net27324);
   U6 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => net27325);
   U7 : INV_X1 port map( A => A, ZN => net27323);
   U1 : OAI21_X1 port map( B1 => net27323, B2 => net27324, A => net27325, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   U3 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U4 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n3);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U3 : XNOR2_X1 port map( A => n6, B => A, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U1 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => n3, B => A, ZN => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n8 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X2 port map( A => n8, B => A, ZN => S);
   U2 : XNOR2_X2 port map( A => B, B => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U7 : CLKBUF_X1 port map( A => A, Z => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6, n8 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => n8, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n6);
   U7 : XNOR2_X1 port map( A => n6, B => A, ZN => S);
   U1 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n6);
   U2 : XNOR2_X1 port map( A => A, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n7 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U4 : INV_X1 port map( A => n7, ZN => n3);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n3, B2 => n2, ZN => Co);
   U1 : CLKBUF_X1 port map( A => A, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n6, n2, n8 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U4 : XNOR2_X1 port map( A => n6, B => n2, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U7 : INV_X1 port map( A => B, ZN => n3);
   U8 : OAI22_X1 port map( A1 => n6, A2 => n8, B1 => n4, B2 => n3, ZN => Co);
   MY_CLK_r_REG588_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n2, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n_1553 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => n6, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => n6, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG624_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1553);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG592_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG622_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   MY_CLK_r_REG613_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG621_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n8, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG665_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n8)
                           ;
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n10 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n10, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG636_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n10
                           );
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_186 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR, clk : in 
         std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n11, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n7, B1 => n2, B2 => n10, ZN => Co);
   MY_CLK_r_REG591_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG669_S1 : DFF_X1 port map( D => Ci_BAR, CK => clk, Q => n7, QN =>
                           n11);
   U3 : XNOR2_X1 port map( A => A, B => n8, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n13, n_1554 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n10, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG590_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1554);
   MY_CLK_r_REG606_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG635_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1555, n_1556 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG670_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1555);
   MY_CLK_r_REG605_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1556);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n3, n_1558 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);
   MY_CLK_r_REG375_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n3, QN => 
                           n_1558);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_204 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => n2, B2 => n1, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n6);
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_205 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n6, B1 => n2, B2 => n1, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n6);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n_1559 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : INV_X1 port map( A => B, ZN => n2);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n2, B2 => n3, A => n1, ZN => Co);
   U5 : FA_X1 port map( A => Ci, B => A, CI => B, CO => n_1559, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n7 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => n7, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_211 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n5, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n5, A2 => n8, B1 => n3, B2 => n2, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : INV_X1 port map( A => Ci, ZN => n2);
   U3 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U5 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U6 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U1 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27478, net27476, n1, n2 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n1, B2 => net27478, A => n2, ZN => Co);
   U2 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => net27476);
   U5 : INV_X1 port map( A => Ci, ZN => net27478);
   U6 : XNOR2_X1 port map( A => net27476, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U4 : INV_X1 port map( A => A, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_216 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n6 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => n3, B2 => n6, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U6 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U4 : INV_X1 port map( A => Ci, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n8 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => n8, ZN => n3);
   U6 : OAI21_X1 port map( B1 => n8, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : CLKBUF_X1 port map( A => B, Z => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_218 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6, n8, n10, n11 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n8, A2 => n10, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n2);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n8);
   U9 : INV_X1 port map( A => B, ZN => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n10);
   U5 : XNOR2_X1 port map( A => A, B => n11, ZN => S);
   U7 : INV_X1 port map( A => A, ZN => n6);
   U8 : XNOR2_X1 port map( A => B, B => Ci, ZN => n11);
   U3 : AND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27497, net27498, net27499, n1, n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U4 : INV_X1 port map( A => B, ZN => net27498);
   U5 : OAI21_X1 port map( B1 => B, B2 => n1, A => Ci, ZN => net27499);
   U6 : INV_X1 port map( A => n1, ZN => net27497);
   U7 : OAI21_X1 port map( B1 => net27497, B2 => net27498, A => net27499, ZN =>
                           Co);
   U1 : CLKBUF_X1 port map( A => A, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27501, net27502, net27503, net27504, n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net27503);
   U4 : INV_X1 port map( A => A, ZN => net27501);
   U5 : INV_X1 port map( A => B, ZN => net27502);
   U6 : INV_X1 port map( A => Ci, ZN => net27504);
   U7 : NAND2_X1 port map( A1 => net27501, A2 => net27502, ZN => n2);
   U8 : NAND2_X1 port map( A1 => net27503, A2 => net27504, ZN => n3);
   U9 : AND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27506, net27507, net27508, n1, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U4 : INV_X1 port map( A => n7, ZN => net27506);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => net27508);
   U6 : INV_X1 port map( A => B, ZN => net27507);
   U8 : OAI21_X1 port map( B1 => net27506, B2 => net27507, A => net27508, ZN =>
                           Co);
   U3 : CLKBUF_X1 port map( A => A, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U8 : INV_X1 port map( A => Ci, ZN => n2);
   U2 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27515, n1, n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => net27515);
   U6 : NAND2_X1 port map( A1 => net27515, A2 => n2, ZN => Co);
   U7 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6, n7, n9, n10 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U5 : INV_X1 port map( A => B, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U1 : NAND2_X1 port map( A1 => n10, A2 => A, ZN => n9);
   U4 : INV_X1 port map( A => n2, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => n10);
   U8 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U10 : NAND2_X1 port map( A1 => n9, A2 => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n9 : std_logic;

begin
   
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n9);
   U2 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U3 : XNOR2_X1 port map( A => A, B => n9, ZN => S);
   U4 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => Ci, B => A, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => n7, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n7, B2 => n6, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U7 : INV_X1 port map( A => n2, ZN => n6);
   U8 : CLKBUF_X1 port map( A => A, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U4 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n4);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => B, ZN => n3);
   U8 : OAI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n6, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n8, ZN => Co);
   MY_CLK_r_REG513_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n7, n8, n10, n11, n12 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => n8, ZN => n4);
   U3 : INV_X1 port map( A => n12, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n11, A2 => n4, B1 => n2, B2 => n10, ZN => Co);
   MY_CLK_r_REG534_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG625_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );
   U4 : BUF_X1 port map( A => A, Z => n12);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n14, ZN => Co)
                           ;
   U3 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   MY_CLK_r_REG535_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG550_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG593_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n14, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG551_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n14
                           );
   MY_CLK_r_REG556_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG623_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1560 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG557_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG564_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1560, QN => 
                           n14);
   MY_CLK_r_REG612_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1561 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG565_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG571_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1561, QN => 
                           n14);
   MY_CLK_r_REG620_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n9, n10, n11, n12, n14, n_1562, n_1563, n_1564 : 
      std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n9, A2 => n14, B1 => n12, B2 => n11, ZN => Co)
                           ;
   MY_CLK_r_REG568_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n12, QN => 
                           n_1562);
   MY_CLK_r_REG586_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n11, QN => 
                           n_1563);
   MY_CLK_r_REG611_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n14);
   MY_CLK_r_REG569_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n9, QN => 
                           n_1564);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n9, n10, n11, n12, n14, n_1565, n_1566, n_1567 : 
      std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n9, A2 => n14, B1 => n12, B2 => n11, ZN => Co)
                           ;
   MY_CLK_r_REG584_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n12, QN => 
                           n_1565);
   MY_CLK_r_REG619_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n11, QN => 
                           n_1566);
   MY_CLK_r_REG638_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n14);
   MY_CLK_r_REG585_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n9, QN => 
                           n_1567);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_271 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR, clk : in 
         std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n2, n_1572 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n2, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U2 : NOR2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   MY_CLK_r_REG583_S1 : DFF_X1 port map( D => B_BAR, CK => clk, Q => n2, QN => 
                           n_1572);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n3, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => n4, ZN => S);
   U2 : NOR2_X1 port map( A1 => n4, A2 => n6, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n4);
   MY_CLK_r_REG582_S1 : DFF_X1 port map( D => B, CK => clk, Q => n3, QN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n8, n9, n12, n_1574 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => n8, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n9, B2 => A, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG581_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG578_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1574);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1575 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG577_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG580_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1575);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n7, n8, n10, n_1576 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n8, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => n7, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U6 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n10, A => n2, ZN => Co);
   MY_CLK_r_REG579_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG573_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1576);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1577 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG574_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG575_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1577);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n_1578 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n6, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => n6, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG602_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1578);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1579 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG603_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG600_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1579);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1580 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG601_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG608_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1580);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1581 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG609_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG598_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1581);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n8, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n11, B1 => n2, B2 => n10, ZN => Co);
   MY_CLK_r_REG599_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG632_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n14, B1 => n12, B2 => n13, ZN => Co)
                           ;
   U3 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   MY_CLK_r_REG528_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG633_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG596_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n14
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n12, n13, n14, n_1582 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U5 : INV_X1 port map( A => n9, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n1, ZN => Co);
   MY_CLK_r_REG560_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1582, QN => 
                           n13);
   MY_CLK_r_REG597_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG630_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n11, B1 => n8, B2 => n1, ZN => Co);
   MY_CLK_r_REG538_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n8, QN => n10
                           );
   MY_CLK_r_REG594_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );
   U3 : XNOR2_X1 port map( A => B, B => n10, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n10, ZN => n4);
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n14, B1 => n12, B2 => n13, ZN => Co)
                           ;
   MY_CLK_r_REG558_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG595_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG628_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n14
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n13, n_1583 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n10, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG552_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1583);
   MY_CLK_r_REG629_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG615_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n14, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG566_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n14
                           );
   MY_CLK_r_REG614_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG627_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_288 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci, clk : in std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component SDFF_X1
      port( D, SI, SE, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n9, n10, n12, n13, n14, n15, n_1584 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n10, B2 => n12, ZN => Co)
                           ;
   MY_CLK_r_REG626_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG649_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   MY_CLK_r_REG572_S1 : SDFF_X1 port map( D => n14, SI => n15, SE => A, CK => 
                           clk, Q => n10, QN => n_1584);
   n14 <= '1';
   n15 <= '0';

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1585, n_1586 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG637_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1585);
   MY_CLK_r_REG589_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1586);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_292 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, n3, n_1588 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => n4, ZN => S);
   MY_CLK_r_REG372_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n3, QN => 
                           n_1588);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_306 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR, clk : in 
         std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n5, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n5, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG374_S1 : DFF_X1 port map( D => Ci_BAR, CK => clk, Q => n5, QN =>
                           n8);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => Ci, B => A, Z => n3);
   U5 : XOR2_X1 port map( A => B, B => n3, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U7 : XNOR2_X1 port map( A => A, B => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U7 : XNOR2_X1 port map( A => n9, B => A, ZN => S);
   U8 : XNOR2_X1 port map( A => B, B => Ci, ZN => n9);
   U1 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U1 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27835, net27836, net27837, n2 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n2);
   U3 : XNOR2_X1 port map( A => n2, B => A, ZN => S);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => net27837);
   U5 : INV_X1 port map( A => B, ZN => net27836);
   U6 : INV_X1 port map( A => A, ZN => net27835);
   U7 : OAI21_X1 port map( B1 => net27835, B2 => net27836, A => net27837, ZN =>
                           Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_317;

architecture SYN_BEHAVIORAL of FA_317 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U7 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U8 : AOI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_318;

architecture SYN_BEHAVIORAL of FA_318 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => A, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => Ci, ZN => n6);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U6 : INV_X1 port map( A => Ci, ZN => n4);
   U7 : INV_X1 port map( A => A, ZN => n3);
   U8 : INV_X1 port map( A => B, ZN => n2);
   U1 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_319;

architecture SYN_BEHAVIORAL of FA_319 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U3 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_320;

architecture SYN_BEHAVIORAL of FA_320 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n8 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U7 : INV_X1 port map( A => A, ZN => n4);
   U8 : INV_X1 port map( A => B, ZN => n3);
   U2 : XNOR2_X1 port map( A => n8, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_321;

architecture SYN_BEHAVIORAL of FA_321 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27856, net27857, net27858, net27859, n1, n2 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => net27858);
   U4 : XNOR2_X1 port map( A => Ci, B => B, ZN => n2);
   U5 : NAND2_X1 port map( A1 => A, A2 => n1, ZN => net27856);
   U6 : INV_X1 port map( A => n1, ZN => net27859);
   U7 : XNOR2_X1 port map( A => n2, B => A, ZN => S);
   U9 : INV_X1 port map( A => Ci, ZN => net27857);
   U8 : AOI22_X1 port map( A1 => net27856, A2 => net27857, B1 => net27858, B2 
                           => net27859, ZN => Co);
   U1 : CLKBUF_X1 port map( A => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_322;

architecture SYN_BEHAVIORAL of FA_322 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U7 : INV_X1 port map( A => Ci, ZN => n1);
   U2 : XNOR2_X1 port map( A => n7, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n7);
   U1 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_323;

architecture SYN_BEHAVIORAL of FA_323 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net35527, net35526, n1 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U5 : AOI21_X1 port map( B1 => A, B2 => Ci, A => B, ZN => net35527);
   U6 : NOR2_X1 port map( A1 => A, A2 => Ci, ZN => net35526);
   U1 : NOR2_X1 port map( A1 => net35527, A2 => net35526, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_324;

architecture SYN_BEHAVIORAL of FA_324 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5, n7, n8, n9, n11 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n2);
   U6 : XNOR2_X1 port map( A => A, B => Ci, ZN => n9);
   U7 : XNOR2_X1 port map( A => n9, B => B, ZN => S);
   U8 : INV_X1 port map( A => A, ZN => n8);
   U9 : INV_X1 port map( A => B, ZN => n7);
   U11 : INV_X1 port map( A => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => n11, A2 => n5, ZN => n3);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n11);
   U1 : AND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_325;

architecture SYN_BEHAVIORAL of FA_325 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net27876, net27877, net27878, net27879, n1 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net27878);
   U4 : INV_X1 port map( A => B, ZN => net27877);
   U6 : INV_X1 port map( A => Ci, ZN => net27879);
   U5 : INV_X1 port map( A => A, ZN => net27876);
   U7 : AOI22_X1 port map( A1 => net27876, A2 => net27877, B1 => net27878, B2 
                           => net27879, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_326;

architecture SYN_BEHAVIORAL of FA_326 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n6 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U1 : XNOR2_X1 port map( A => A, B => n6, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_327;

architecture SYN_BEHAVIORAL of FA_327 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n8 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => n8);
   U8 : XNOR2_X1 port map( A => n8, B => A, ZN => S);
   U2 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_328;

architecture SYN_BEHAVIORAL of FA_328 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U4 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_329;

architecture SYN_BEHAVIORAL of FA_329 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n7, n10 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n7, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n10, ZN => Co);
   MY_CLK_r_REG412_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n10)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_330;

architecture SYN_BEHAVIORAL of FA_330 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n_1589 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n4);
   U3 : INV_X1 port map( A => B, ZN => n3);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U6 : FA_X1 port map( A => A, B => B, CI => Ci, CO => n_1589, S => S);
   U1 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_331;

architecture SYN_BEHAVIORAL of FA_331 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_332;

architecture SYN_BEHAVIORAL of FA_332 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_333;

architecture SYN_BEHAVIORAL of FA_333 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n8, n_1590 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => n6, B => B, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n6, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   MY_CLK_r_REG529_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1590);
   U7 : INV_X1 port map( A => n3, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_334;

architecture SYN_BEHAVIORAL of FA_334 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n6, n7, n9, n_1591, n_1592 : std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n6, B => n7, Z => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => n7, A => n6, ZN => n3);
   MY_CLK_r_REG471_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => 
                           n_1591);
   MY_CLK_r_REG561_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1592);
   U1 : XNOR2_X1 port map( A => n1, B => n9, ZN => S);
   U6 : INV_X1 port map( A => A, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_335;

architecture SYN_BEHAVIORAL of FA_335 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1593 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG483_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG539_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1593);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_336;

architecture SYN_BEHAVIORAL of FA_336 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n7, n8, n9, n11, n_1594, n_1595, n_1596 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n3);
   MY_CLK_r_REG484_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1594);
   MY_CLK_r_REG498_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1595);
   MY_CLK_r_REG559_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1596);
   U1 : XNOR2_X1 port map( A => n9, B => n8, ZN => n11);
   U2 : XNOR2_X1 port map( A => n11, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_337;

architecture SYN_BEHAVIORAL of FA_337 is

   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n8, n9, n10, n12, n13, n14, n15 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U3 : INV_X1 port map( A => n10, ZN => n2);
   U5 : INV_X1 port map( A => n9, ZN => n1);
   MY_CLK_r_REG499_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n14
                           );
   MY_CLK_r_REG504_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n15)
                           ;
   MY_CLK_r_REG553_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : CLKBUF_X1 port map( A => n4, Z => n13);
   U4 : XNOR2_X1 port map( A => n14, B => n15, ZN => n4);
   U6 : OAI22_X2 port map( A1 => n13, A2 => n12, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_338;

architecture SYN_BEHAVIORAL of FA_338 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U3 : INV_X1 port map( A => n10, ZN => n2);
   U5 : INV_X1 port map( A => n9, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG505_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG511_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG567_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_339;

architecture SYN_BEHAVIORAL of FA_339 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6, n7, n_1597, n_1598 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U5 : XOR2_X1 port map( A => B, B => Ci, Z => n4);
   U6 : XOR2_X1 port map( A => n7, B => n6, Z => S);
   MY_CLK_r_REG512_S1 : DFF_X1 port map( D => A, CK => clk, Q => n7, QN => 
                           n_1597);
   MY_CLK_r_REG526_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n6, QN => 
                           n_1598);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_340;

architecture SYN_BEHAVIORAL of FA_340 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U3 : INV_X1 port map( A => n10, ZN => n2);
   U5 : INV_X1 port map( A => n9, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n12, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG527_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG533_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG587_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_342;

architecture SYN_BEHAVIORAL of FA_342 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_366;

architecture SYN_BEHAVIORAL of FA_366 is

begin
   S <= B;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_368;

architecture SYN_BEHAVIORAL of FA_368 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);
   U2 : AND2_X1 port map( A1 => A, A2 => B, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_369;

architecture SYN_BEHAVIORAL of FA_369 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U4 : INV_X1 port map( A => B, ZN => n2);
   U2 : NOR2_X1 port map( A1 => n4, A2 => n2, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U1 : XNOR2_X1 port map( A => n2, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_370;

architecture SYN_BEHAVIORAL of FA_370 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U1 : NOR2_X1 port map( A1 => n3, A2 => n5, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_371;

architecture SYN_BEHAVIORAL of FA_371 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1605, n_1606 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   MY_CLK_r_REG610_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1605);
   MY_CLK_r_REG576_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n7, QN => 
                           n_1606);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_372;

architecture SYN_BEHAVIORAL of FA_372 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U4 : INV_X1 port map( A => B, ZN => n2);
   U2 : NOR2_X1 port map( A1 => n4, A2 => n2, ZN => Co);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U1 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_373;

architecture SYN_BEHAVIORAL of FA_373 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_374;

architecture SYN_BEHAVIORAL of FA_374 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_378 is

   port( A, B : in std_logic;  S, Co : out std_logic;  clk, Ci : in std_logic);

end FA_378;

architecture SYN_BEHAVIORAL of FA_378 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n7, n8, n10, n_1608, n_1609 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n10, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG641_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1608);
   MY_CLK_r_REG631_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1609);
   U4 : INV_X1 port map( A => Ci, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_387;

architecture SYN_BEHAVIORAL of FA_387 is

begin
   S <= A;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_388 is

   port( A, Ci : in std_logic;  Co : out std_logic;  B_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_388;

architecture SYN_BEHAVIORAL of FA_388 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n6 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U1 : INV_X1 port map( A => B_BAR, ZN => n6);
   U4 : NOR2_X1 port map( A1 => n2, A2 => B_BAR, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => n6, ZN => S_BAR);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_389 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR, clk : in 
         std_logic);

end FA_389;

architecture SYN_BEHAVIORAL of FA_389 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n13, n_1614 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n12, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n13, B1 => n10, B2 => n9, ZN => Co);
   MY_CLK_r_REG365_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1614);
   MY_CLK_r_REG440_S1 : DFF_X1 port map( D => B_BAR, CK => clk, Q => n9, QN => 
                           n12);
   MY_CLK_r_REG427_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_390 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR, clk : in 
         std_logic);

end FA_390;

architecture SYN_BEHAVIORAL of FA_390 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n_1615, n_1616 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n9, ZN => Co);
   MY_CLK_r_REG643_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1615);
   MY_CLK_r_REG426_S1 : DFF_X1 port map( D => B_BAR, CK => clk, Q => n9, QN => 
                           n_1616);
   MY_CLK_r_REG370_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XNOR2_X1 port map( A => n10, B => n9, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_391;

architecture SYN_BEHAVIORAL of FA_391 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1617, n_1618 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n14, B2 => n13, ZN => Co)
                           ;
   MY_CLK_r_REG357_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1617, QN => 
                           n14);
   MY_CLK_r_REG371_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1618, QN => 
                           n13);
   MY_CLK_r_REG424_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_392;

architecture SYN_BEHAVIORAL of FA_392 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1619, n_1620 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n14, B2 => n13, ZN => Co)
                           ;
   MY_CLK_r_REG363_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1619, QN => 
                           n14);
   MY_CLK_r_REG425_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1620, QN => 
                           n13);
   MY_CLK_r_REG438_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_393;

architecture SYN_BEHAVIORAL of FA_393 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n8, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => n7, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n11, B1 => n2, B2 => n10, ZN => Co);
   MY_CLK_r_REG439_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG449_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_394;

architecture SYN_BEHAVIORAL of FA_394 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n_1621, n_1622, n_1623 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n3);
   U5 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n2);
   MY_CLK_r_REG336_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1621);
   MY_CLK_r_REG450_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1622);
   MY_CLK_r_REG453_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1623);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_395;

architecture SYN_BEHAVIORAL of FA_395 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1624 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG454_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG462_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1624);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_396;

architecture SYN_BEHAVIORAL of FA_396 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n8, n10, n_1625 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n8, B2 => A, A => n7, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n10, A => n1, ZN => Co);
   MY_CLK_r_REG463_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG489_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1625);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_397;

architecture SYN_BEHAVIORAL of FA_397 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6, n7, n_1626, n_1627 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n1);
   U3 : OAI21_X1 port map( B1 => n7, B2 => A, A => n6, ZN => n2);
   U4 : XOR2_X1 port map( A => n6, B => n7, Z => n3);
   U5 : XOR2_X1 port map( A => A, B => n3, Z => S);
   MY_CLK_r_REG490_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => 
                           n_1626);
   MY_CLK_r_REG477_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1627);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_398;

architecture SYN_BEHAVIORAL of FA_398 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28155, net28157, n1, n5, n6, n8, n_1628 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n5, ZN => n1);
   U2 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U3 : OAI21_X1 port map( B1 => A, B2 => n6, A => n5, ZN => net28157);
   U5 : INV_X1 port map( A => A, ZN => net28155);
   U6 : OAI21_X1 port map( B1 => net28155, B2 => n8, A => net28157, ZN => Co);
   MY_CLK_r_REG478_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => n8);
   MY_CLK_r_REG480_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n5, QN => 
                           n_1628);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_399;

architecture SYN_BEHAVIORAL of FA_399 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6, n_1629 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => n6, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG486_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1629);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_400;

architecture SYN_BEHAVIORAL of FA_400 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n8, n9, n11, n_1630 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => n8, ZN => S);
   U3 : XNOR2_X1 port map( A => n9, B => A, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U6 : OAI21_X1 port map( B1 => n9, B2 => A, A => n8, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n11, A => n2, ZN => Co);
   MY_CLK_r_REG487_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n11)
                           ;
   MY_CLK_r_REG503_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1630);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_401;

architecture SYN_BEHAVIORAL of FA_401 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n5, n_1631 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : OAI21_X1 port map( B1 => A, B2 => B, A => n5, ZN => n2);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n1);
   MY_CLK_r_REG509_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n5, QN => 
                           n_1631);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_402;

architecture SYN_BEHAVIORAL of FA_402 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5, n6, n8, n9, n11, n12 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => n6, ZN => S);
   U3 : XNOR2_X1 port map( A => n9, B => n8, ZN => n6);
   U4 : NAND2_X1 port map( A1 => n9, A2 => A, ZN => n5);
   U6 : INV_X1 port map( A => A, ZN => n3);
   U8 : AOI22_X1 port map( A1 => n5, A2 => n12, B1 => n3, B2 => n11, ZN => Co);
   MY_CLK_r_REG510_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n11)
                           ;
   MY_CLK_r_REG524_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_403;

architecture SYN_BEHAVIORAL of FA_403 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n9, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n13, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG306_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG525_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG531_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n14
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_404;

architecture SYN_BEHAVIORAL of FA_404 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n_1632, n_1633, n_1634 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n1);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n2);
   MY_CLK_r_REG417_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1632);
   MY_CLK_r_REG532_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1633);
   MY_CLK_r_REG522_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1634);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_405;

architecture SYN_BEHAVIORAL of FA_405 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n10, ZN => S);
   U4 : INV_X1 port map( A => n9, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n10, B2 => n9, A => n8, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n3, A => n2, ZN => Co);
   MY_CLK_r_REG428_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG523_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG548_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_406;

architecture SYN_BEHAVIORAL of FA_406 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1635, n_1636 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG445_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1635, QN => 
                           n13);
   MY_CLK_r_REG549_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1636, QN => 
                           n14);
   MY_CLK_r_REG520_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_407;

architecture SYN_BEHAVIORAL of FA_407 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1637 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n8, B => n10, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n13, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG495_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG521_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG546_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1637);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_408;

architecture SYN_BEHAVIORAL of FA_408 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1638 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n9, B => n8, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n13, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG451_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG547_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG516_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1638);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_409;

architecture SYN_BEHAVIORAL of FA_409 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n11, n12, n_1639 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => n8, B => n3, ZN => S);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n1);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n2);
   MY_CLK_r_REG492_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG517_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1639);
   MY_CLK_r_REG544_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );
   U1 : XNOR2_X1 port map( A => n11, B => n12, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_410;

architecture SYN_BEHAVIORAL of FA_410 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n7, n8, n9, n10, n12, n13, n_1640 : std_logic;

begin
   
   U6 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n13, B2 => n12, A => n2, ZN => Co);
   U2 : XNOR2_X1 port map( A => n8, B => n10, ZN => n7);
   MY_CLK_r_REG481_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG545_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG540_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1640);
   U1 : XNOR2_X1 port map( A => n7, B => n9, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_411;

architecture SYN_BEHAVIORAL of FA_411 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1641 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n9, B => n8, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n1, ZN => Co);
   MY_CLK_r_REG491_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG541_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG542_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1641);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_412;

architecture SYN_BEHAVIORAL of FA_412 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n5, n8, n9, n10, n12, n15, n_1642 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n9, B => n5, ZN => S);
   U3 : XNOR2_X1 port map( A => n10, B => n8, ZN => n5);
   U6 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n15, B2 => n12, A => n2, ZN => Co);
   MY_CLK_r_REG496_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n15
                           );
   MY_CLK_r_REG543_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG555_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1642);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_413;

architecture SYN_BEHAVIORAL of FA_413 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n9, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n14, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG506_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n14
                           );
   MY_CLK_r_REG554_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG562_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_414;

architecture SYN_BEHAVIORAL of FA_414 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1643, n_1644 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG519_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1643, QN => 
                           n13);
   MY_CLK_r_REG563_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1644, QN => 
                           n14);
   MY_CLK_r_REG607_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_415;

architecture SYN_BEHAVIORAL of FA_415 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n6, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U7 : XNOR2_X1 port map( A => A, B => B, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_420;

architecture SYN_BEHAVIORAL of FA_420 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : XOR2_X1 port map( A => n3, B => B, Z => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n4);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : OAI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_429;

architecture SYN_BEHAVIORAL of FA_429 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n6, n10, n11, n_1646, n_1647, n_1648 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   MY_CLK_r_REG642_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n_1646, QN =>
                           n10);
   MY_CLK_r_REG645_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1647, QN => 
                           n11);
   MY_CLK_r_REG377_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1648);
   U3 : XOR2_X1 port map( A => n10, B => n11, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_430;

architecture SYN_BEHAVIORAL of FA_430 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n10, n12, n13, n14, n_1649 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG646_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n13);
   MY_CLK_r_REG647_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1649, QN => 
                           n14);
   MY_CLK_r_REG373_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XOR2_X1 port map( A => n13, B => n14, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_431;

architecture SYN_BEHAVIORAL of FA_431 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n8, n12, n13, n14, n_1650, n_1651 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n13, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG648_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1650, QN => 
                           n13);
   MY_CLK_r_REG650_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1651, QN => 
                           n14);
   MY_CLK_r_REG376_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );
   U3 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_432;

architecture SYN_BEHAVIORAL of FA_432 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n8, n9, n10, n12, n14, n_1652 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n10, B => n9, Z => n4);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n12, B1 => n10, B2 => n14, ZN => Co)
                           ;
   MY_CLK_r_REG651_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1652);
   MY_CLK_r_REG658_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG369_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n12
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_433;

architecture SYN_BEHAVIORAL of FA_433 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n9, n13, n14, n15, n_1653, n_1654 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n9, ZN => S);
   U6 : OAI22_X1 port map( A1 => n15, A2 => n14, B1 => n4, B2 => n13, ZN => Co)
                           ;
   MY_CLK_r_REG659_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1653, QN => 
                           n15);
   MY_CLK_r_REG656_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1654, QN => 
                           n14);
   MY_CLK_r_REG644_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => n13
                           );
   U4 : XNOR2_X1 port map( A => n14, B => n15, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_434;

architecture SYN_BEHAVIORAL of FA_434 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n4, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n14, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG657_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n14
                           );
   MY_CLK_r_REG652_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG362_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   U2 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_435;

architecture SYN_BEHAVIORAL of FA_435 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1655 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n8, B => n9, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n1, ZN => Co);
   MY_CLK_r_REG653_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG655_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG364_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1655);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_436;

architecture SYN_BEHAVIORAL of FA_436 is

   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n_1656 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : INV_X1 port map( A => B, ZN => n2);
   U3 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U5 : FA_X1 port map( A => B, B => A, CI => Ci, CO => n_1656, S => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_437;

architecture SYN_BEHAVIORAL of FA_437 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n8, n9, n11, n_1657 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => A, B => n8, ZN => n5);
   U3 : XNOR2_X1 port map( A => n5, B => n9, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U6 : OAI21_X1 port map( B1 => n9, B2 => A, A => n8, ZN => n2);
   MY_CLK_r_REG343_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n11)
                           ;
   MY_CLK_r_REG341_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1657);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n11, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_438;

architecture SYN_BEHAVIORAL of FA_438 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_439;

architecture SYN_BEHAVIORAL of FA_439 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n7, n8, n10, n11 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n8, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n7, B2 => n8, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n10, B2 => n11, A => n1, ZN => Co);
   MY_CLK_r_REG345_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n10)
                           ;
   MY_CLK_r_REG334_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n11)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_440;

architecture SYN_BEHAVIORAL of FA_440 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n11, n12 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n9, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => n8, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n11, B2 => n12, A => n1, ZN => Co);
   MY_CLK_r_REG335_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => n11)
                           ;
   MY_CLK_r_REG663_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n12)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_441;

architecture SYN_BEHAVIORAL of FA_441 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n7, n9 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n7, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U5 : OAI21_X1 port map( B1 => n7, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n9, A => n1, ZN => Co);
   MY_CLK_r_REG323_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_442;

architecture SYN_BEHAVIORAL of FA_442 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U5 : INV_X1 port map( A => Ci, ZN => n2);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U1 : AOI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_443;

architecture SYN_BEHAVIORAL of FA_443 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n7, n9 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => n7, ZN => n5);
   U3 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n9, ZN => Co);
   MY_CLK_r_REG313_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_444;

architecture SYN_BEHAVIORAL of FA_444 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_445;

architecture SYN_BEHAVIORAL of FA_445 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28326, net28327, n1, n6, n7, n9, n10 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => net28326, A2 => net28327, B1 => n10, B2 => n9,
                           ZN => Co);
   U2 : XNOR2_X1 port map( A => n1, B => n6, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => n7, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => net28326);
   U6 : INV_X1 port map( A => Ci, ZN => net28327);
   MY_CLK_r_REG317_S1 : DFF_X1 port map( D => A, CK => clk, Q => n7, QN => n10)
                           ;
   MY_CLK_r_REG303_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_446;

architecture SYN_BEHAVIORAL of FA_446 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6, n7, n_1658, n_1659 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : NOR2_X1 port map( A1 => n6, A2 => n7, ZN => n1);
   U3 : AOI21_X1 port map( B1 => n7, B2 => n6, A => Ci, ZN => n2);
   U4 : XNOR2_X1 port map( A => n3, B => n6, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => n7, ZN => n3);
   MY_CLK_r_REG304_S1 : DFF_X1 port map( D => A, CK => clk, Q => n7, QN => 
                           n_1658);
   MY_CLK_r_REG296_S1 : DFF_X1 port map( D => B, CK => clk, Q => n6, QN => 
                           n_1659);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_447;

architecture SYN_BEHAVIORAL of FA_447 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28334, net28335, n1, n6, n7, n8, n10, n11, n12 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n7, ZN => S);
   U5 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => net28334);
   U7 : INV_X1 port map( A => n6, ZN => net28335);
   MY_CLK_r_REG295_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n11)
                           ;
   MY_CLK_r_REG290_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n10)
                           ;
   MY_CLK_r_REG416_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => n12
                           );
   U2 : AOI22_X1 port map( A1 => net28334, A2 => net28335, B1 => n11, B2 => n10
                           , ZN => Co);
   U3 : XNOR2_X1 port map( A => n11, B => n12, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_448;

architecture SYN_BEHAVIORAL of FA_448 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n6, n10, n12, n13, n_1660 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : NAND2_X1 port map( A1 => n10, A2 => B, ZN => n3);
   U2 : AOI22_X1 port map( A1 => n12, A2 => n4, B1 => n3, B2 => n13, ZN => Co);
   MY_CLK_r_REG294_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG429_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n_1660, QN =>
                           n13);
   U1 : XNOR2_X1 port map( A => n12, B => n13, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_449;

architecture SYN_BEHAVIORAL of FA_449 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28348, net33793, n1, n2, n6, n7, n8, n10, n11, n_1661 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => n8, B => n6, ZN => n1);
   U5 : AND2_X1 port map( A1 => n11, A2 => n6, ZN => net28348);
   U6 : AND2_X1 port map( A1 => n6, A2 => n10, ZN => net33793);
   U7 : XNOR2_X1 port map( A => net33793, B => net28348, ZN => n2);
   U8 : OAI21_X1 port map( B1 => n11, B2 => n10, A => n2, ZN => Co);
   MY_CLK_r_REG287_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => n11)
                           ;
   MY_CLK_r_REG288_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => n10)
                           ;
   MY_CLK_r_REG446_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n6, QN => 
                           n_1661);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_450;

architecture SYN_BEHAVIORAL of FA_450 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n5, n8, n9, n11, n12 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => n9, B => n8, ZN => n5);
   U6 : OAI21_X1 port map( B1 => n9, B2 => n8, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n12, B2 => n11, A => n2, ZN => Co);
   MY_CLK_r_REG289_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG276_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n11)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_451;

architecture SYN_BEHAVIORAL of FA_451 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n7, n8, n9, n_1662, n_1663, n_1664 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n2, B => n8, ZN => S);
   U4 : XNOR2_X1 port map( A => n9, B => n7, ZN => n2);
   U5 : AOI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n4);
   U6 : NOR2_X1 port map( A1 => n9, A2 => n8, ZN => n3);
   U1 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => Co);
   MY_CLK_r_REG279_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1662);
   MY_CLK_r_REG272_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1663);
   MY_CLK_r_REG452_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1664);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_452;

architecture SYN_BEHAVIORAL of FA_452 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n14 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n10, ZN => S);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   MY_CLK_r_REG275_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG200_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n14)
                           ;
   MY_CLK_r_REG493_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => n13
                           );
   U2 : OAI21_X1 port map( B1 => n12, B2 => n14, A => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => n13, B => n14, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_453;

architecture SYN_BEHAVIORAL of FA_453 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n10, n11, n12, n14, n15, n_1665, n_1666 : std_logic;

begin
   
   U3 : OAI21_X1 port map( B1 => n11, B2 => n12, A => n10, ZN => n1);
   U4 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n1, ZN => Co);
   U5 : FA_X1 port map( A => n12, B => n11, CI => n10, CO => n_1665, S => S);
   MY_CLK_r_REG268_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n14
                           );
   MY_CLK_r_REG410_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n15
                           );
   MY_CLK_r_REG482_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n_1666);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_454;

architecture SYN_BEHAVIORAL of FA_454 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1667, n_1668 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n8, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG411_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => 
                           n_1667);
   MY_CLK_r_REG432_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1668);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_455;

architecture SYN_BEHAVIORAL of FA_455 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n_1669, n_1670, n_1671 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => n9, B => n7, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n1);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n2);
   MY_CLK_r_REG433_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1669);
   MY_CLK_r_REG441_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1670);
   MY_CLK_r_REG497_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1671);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_456;

architecture SYN_BEHAVIORAL of FA_456 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n11, n12, n_1672 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => n8, ZN => S);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n1);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n2);
   MY_CLK_r_REG442_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG457_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1672);
   MY_CLK_r_REG507_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );
   U2 : XNOR2_X1 port map( A => n11, B => n12, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_457;

architecture SYN_BEHAVIORAL of FA_457 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n5, n6, n7, n8, n12, n13, n14, n15, n17, n18, n_1673, n_1674 : 
      std_logic;

begin
   
   U2 : XOR2_X1 port map( A => n15, B => n12, Z => S);
   U3 : XOR2_X1 port map( A => B, B => Ci, Z => n2);
   U4 : NAND2_X1 port map( A1 => n13, A2 => n18, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => Co);
   U7 : NAND2_X1 port map( A1 => n15, A2 => n14, ZN => n7);
   U8 : XNOR2_X1 port map( A => n6, B => n5, ZN => n8);
   U9 : NAND2_X1 port map( A1 => n13, A2 => n17, ZN => n5);
   MY_CLK_r_REG458_S1 : DFF_X1 port map( D => A, CK => clk, Q => n15, QN => n18
                           );
   MY_CLK_r_REG464_S1 : DFF_X1 port map( D => B, CK => clk, Q => n14, QN => n17
                           );
   MY_CLK_r_REG518_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n13, QN => 
                           n_1673);
   MY_CLK_r_REG465_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n12, QN => 
                           n_1674);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_458;

architecture SYN_BEHAVIORAL of FA_458 is

   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n10, n13, n14, n16, n17, n_1675, n_1676, n_1677, 
      n_1678, n_1679 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   MY_CLK_r_REG467_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n14, QN => 
                           n_1675);
   MY_CLK_r_REG475_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n13, QN => 
                           n_1676);
   MY_CLK_r_REG466_S1 : DFF_X1 port map( D => A, CK => clk, Q => n_1677, QN => 
                           n16);
   MY_CLK_r_REG476_S1 : DFF_X1 port map( D => n1, CK => clk, Q => n_1678, QN =>
                           n17);
   MY_CLK_r_REG468_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n10, QN => 
                           n_1679);
   U2 : XNOR2_X1 port map( A => n16, B => n17, ZN => S);
   U1 : OAI21_X2 port map( B1 => n14, B2 => n13, A => n10, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_459;

architecture SYN_BEHAVIORAL of FA_459 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6, n7, n_1680, n_1681 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   MY_CLK_r_REG485_S1 : DFF_X1 port map( D => B, CK => clk, Q => n7, QN => 
                           n_1680);
   MY_CLK_r_REG472_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n6, QN => 
                           n_1681);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_461;

architecture SYN_BEHAVIORAL of FA_461 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_463;

architecture SYN_BEHAVIORAL of FA_463 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U1 : XNOR2_X1 port map( A => n5, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_464;

architecture SYN_BEHAVIORAL of FA_464 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_19 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_19;

architecture SYN_rtl of HA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_479 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic);

end FA_479;

architecture SYN_BEHAVIORAL of FA_479 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : NOR2_X1 port map( A1 => n4, A2 => B_BAR, ZN => Co);
   U3 : INV_X1 port map( A => B_BAR, ZN => n6);
   U4 : INV_X1 port map( A => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_480 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic);

end FA_480;

architecture SYN_BEHAVIORAL of FA_480 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => A_BAR, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_482 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic);

end FA_482;

architecture SYN_BEHAVIORAL of FA_482 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U2 : NOR2_X1 port map( A1 => n4, A2 => B_BAR, ZN => Co);
   U3 : INV_X1 port map( A => B_BAR, ZN => n6);
   U4 : INV_X1 port map( A => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_483;

architecture SYN_BEHAVIORAL of FA_483 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_484;

architecture SYN_BEHAVIORAL of FA_484 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n2, B2 => n3, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_24 is

   port( B : in std_logic;  C, S_BAR : out std_logic;  A_BAR : in std_logic);

end HA_24;

architecture SYN_rtl of HA_24 is

begin
   S_BAR <= A_BAR;

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_485 is

   port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_485;

architecture SYN_BEHAVIORAL of FA_485 is

begin
   S_BAR <= A_BAR;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_486 is

   port( A, Ci : in std_logic;  Co : out std_logic;  B_BAR : in std_logic;  
         S_BAR : out std_logic);

end FA_486;

architecture SYN_BEHAVIORAL of FA_486 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n6 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => n6, Z => S_BAR);
   U1 : NOR2_X1 port map( A1 => n2, A2 => B_BAR, ZN => Co);
   U4 : INV_X1 port map( A => B_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_488 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_488;

architecture SYN_BEHAVIORAL of FA_488 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_492 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_492;

architecture SYN_BEHAVIORAL of FA_492 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n6, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_493 is

   port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic);

end FA_493;

architecture SYN_BEHAVIORAL of FA_493 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => n6, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => Ci_BAR, B1 => n2, B2 => n1, ZN => Co
                           );
   U4 : INV_X1 port map( A => Ci_BAR, ZN => n6);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_494;

architecture SYN_BEHAVIORAL of FA_494 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28552, net28553, n1, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U2 : XNOR2_X1 port map( A => n1, B => B, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => net28552);
   U5 : INV_X1 port map( A => B, ZN => net28553);
   U3 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n4);
   U6 : OAI21_X1 port map( B1 => net28552, B2 => net28553, A => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_495;

architecture SYN_BEHAVIORAL of FA_495 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6, n7, n_1693, n_1694 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);
   MY_CLK_r_REG488_S1 : DFF_X1 port map( D => n5, CK => clk, Q => n6, QN => 
                           n_1693);
   MY_CLK_r_REG479_S1 : DFF_X2 port map( D => A, CK => clk, Q => n7, QN => 
                           n_1694);
   U2 : XNOR2_X1 port map( A => n7, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_496;

architecture SYN_BEHAVIORAL of FA_496 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n8 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => n8, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_497;

architecture SYN_BEHAVIORAL of FA_497 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n7, n6, n8, n_1695, n_1696 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => B, B => Ci, ZN => n7);
   MY_CLK_r_REG502_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => 
                           n_1695);
   MY_CLK_r_REG508_S1 : DFF_X1 port map( D => n7, CK => clk, Q => n6, QN => 
                           n_1696);
   U2 : XNOR2_X1 port map( A => n8, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_498;

architecture SYN_BEHAVIORAL of FA_498 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_499;

architecture SYN_BEHAVIORAL of FA_499 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_500;

architecture SYN_BEHAVIORAL of FA_500 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n5 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n3);
   U1 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_501;

architecture SYN_BEHAVIORAL of FA_501 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => n7, B => A, ZN => S);
   U7 : XNOR2_X1 port map( A => Ci, B => B, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_502;

architecture SYN_BEHAVIORAL of FA_502 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_503;

architecture SYN_BEHAVIORAL of FA_503 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_506;

architecture SYN_BEHAVIORAL of FA_506 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_507;

architecture SYN_BEHAVIORAL of FA_507 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_508;

architecture SYN_BEHAVIORAL of FA_508 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_26 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_26;

architecture SYN_rtl of HA_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n1);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_509;

architecture SYN_BEHAVIORAL of FA_509 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_511;

architecture SYN_BEHAVIORAL of FA_511 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_515 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_515;

architecture SYN_BEHAVIORAL of FA_515 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_516 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_516;

architecture SYN_BEHAVIORAL of FA_516 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n13, n14, n_1698 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => n9, ZN => S);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n2);
   U5 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n3);
   MY_CLK_r_REG355_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1698);
   MY_CLK_r_REG347_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n14)
                           ;
   MY_CLK_r_REG423_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n13
                           );
   U6 : XNOR2_X1 port map( A => n13, B => n14, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_517 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_517;

architecture SYN_BEHAVIORAL of FA_517 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_518 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_518;

architecture SYN_BEHAVIORAL of FA_518 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4, n5, n9, n10, n11, n13, n14, n_1699 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => n9, ZN => S);
   U4 : INV_X1 port map( A => n11, ZN => n4);
   U6 : OAI21_X1 port map( B1 => n11, B2 => n10, A => n9, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n13, A => n2, ZN => Co);
   MY_CLK_r_REG346_S1 : DFF_X1 port map( D => A, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG422_S1 : DFF_X1 port map( D => B, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG436_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => 
                           n_1699);
   U1 : XNOR2_X1 port map( A => n13, B => n14, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_519 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_519;

architecture SYN_BEHAVIORAL of FA_519 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4, n8, n9, n10, n12, n13, n_1700 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n10, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n9, B => n8, ZN => n4);
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n1, ZN => Co);
   MY_CLK_r_REG331_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n12
                           );
   MY_CLK_r_REG437_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n13)
                           ;
   MY_CLK_r_REG420_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1700);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_520 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_520;

architecture SYN_BEHAVIORAL of FA_520 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n5, n10, n11, n12, n14, n15, n16 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => n12, ZN => S);
   U6 : OAI21_X1 port map( B1 => n11, B2 => n12, A => n10, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n2, ZN => Co);
   MY_CLK_r_REG661_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n14
                           );
   MY_CLK_r_REG421_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n15
                           );
   MY_CLK_r_REG327_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n16);
   U1 : XNOR2_X1 port map( A => n15, B => n16, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_521 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_521;

architecture SYN_BEHAVIORAL of FA_521 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n9, n10, n11, n12, n14, n15, n16 : std_logic;

begin
   
   U6 : OAI21_X1 port map( B1 => n11, B2 => n12, A => n10, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n15, B2 => n14, A => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => n9, B => n11, ZN => S);
   MY_CLK_r_REG318_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n15
                           );
   MY_CLK_r_REG330_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n14
                           );
   MY_CLK_r_REG418_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n10, QN => 
                           n16);
   U1 : XNOR2_X1 port map( A => n15, B => n16, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_522 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_522;

architecture SYN_BEHAVIORAL of FA_522 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n7, n8, n9, n10, n12, n13, n_1701 : std_logic;

begin
   
   U5 : OAI21_X1 port map( B1 => n9, B2 => n10, A => n8, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n13, B2 => n12, A => n1, ZN => Co);
   U1 : XNOR2_X1 port map( A => n8, B => n10, ZN => n7);
   U2 : XNOR2_X1 port map( A => n7, B => n9, ZN => S);
   MY_CLK_r_REG325_S1 : DFF_X1 port map( D => A, CK => clk, Q => n10, QN => n13
                           );
   MY_CLK_r_REG419_S1 : DFF_X1 port map( D => B, CK => clk, Q => n9, QN => n12)
                           ;
   MY_CLK_r_REG430_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1701);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_523 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_523;

architecture SYN_BEHAVIORAL of FA_523 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7, n8, n9, n_1702, n_1703, n_1704 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => n9, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n3);
   U5 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n2);
   MY_CLK_r_REG307_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1702);
   MY_CLK_r_REG431_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => 
                           n_1703);
   MY_CLK_r_REG447_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => 
                           n_1704);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_524 is

   port( A, B : in std_logic;  S, Co : out std_logic;  clk, Ci_BAR : in 
         std_logic);

end FA_524;

architecture SYN_BEHAVIORAL of FA_524 is

   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n10, n11, n12, n13, n15, n16, n_1705, n_1706 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n11, B => n10, ZN => S);
   U5 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => n6);
   MY_CLK_r_REG455_S1 : DFF_X1 port map( D => Ci_BAR, CK => clk, Q => n13, QN 
                           => n_1705);
   MY_CLK_r_REG314_S1 : DFF_X1 port map( D => A, CK => clk, Q => n12, QN => n15
                           );
   MY_CLK_r_REG448_S1 : DFF_X1 port map( D => B, CK => clk, Q => n11, QN => n16
                           );
   MY_CLK_r_REG315_S1 : DFF_X1 port map( D => n7, CK => clk, Q => n10, QN => 
                           n_1706);
   U2 : XOR2_X1 port map( A => Ci_BAR, B => A, Z => n7);
   U1 : AOI22_X2 port map( A1 => n6, A2 => n13, B1 => n15, B2 => n16, ZN => Co)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_525 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_525;

architecture SYN_BEHAVIORAL of FA_525 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n5, n6, n7, n12, n13, n14, n16, n17, n18, n_1707, n_1708 : 
      std_logic;

begin
   
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n7);
   U5 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => n6);
   U6 : INV_X1 port map( A => Ci, ZN => n5);
   U8 : INV_X1 port map( A => n12, ZN => n3);
   U9 : AOI22_X1 port map( A1 => n6, A2 => n14, B1 => n16, B2 => n3, ZN => Co);
   MY_CLK_r_REG469_S1 : DFF_X1 port map( D => n5, CK => clk, Q => n14, QN => 
                           n_1707);
   MY_CLK_r_REG300_S1 : DFF_X1 port map( D => A, CK => clk, Q => n13, QN => n16
                           );
   MY_CLK_r_REG456_S1 : DFF_X1 port map( D => B, CK => clk, Q => n12, QN => n18
                           );
   MY_CLK_r_REG301_S1 : DFF_X1 port map( D => n7, CK => clk, Q => n_1708, QN =>
                           n17);
   U1 : XNOR2_X1 port map( A => n17, B => n18, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_526 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_526;

architecture SYN_BEHAVIORAL of FA_526 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n10, n11, n_1709, n_1710 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => Co);
   MY_CLK_r_REG470_S1 : DFF_X1 port map( D => B, CK => clk, Q => n_1709, QN => 
                           n11);
   MY_CLK_r_REG305_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n_1710, QN =>
                           n10);
   U1 : XNOR2_X1 port map( A => n10, B => n11, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_527 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_527;

architecture SYN_BEHAVIORAL of FA_527 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => B, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => Ci, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_528 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_528;

architecture SYN_BEHAVIORAL of FA_528 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n7 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U1 : XNOR2_X1 port map( A => B, B => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_530 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_530;

architecture SYN_BEHAVIORAL of FA_530 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6, n8, n9, n_1711, n_1712 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n8, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   MY_CLK_r_REG530_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n9, QN => 
                           n_1711);
   MY_CLK_r_REG494_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n8, QN => 
                           n_1712);
   U3 : XNOR2_X1 port map( A => n2, B => n6, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n6);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_531 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_531;

architecture SYN_BEHAVIORAL of FA_531 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_532 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_532;

architecture SYN_BEHAVIORAL of FA_532 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_533 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_533;

architecture SYN_BEHAVIORAL of FA_533 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_534 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_534;

architecture SYN_BEHAVIORAL of FA_534 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_535 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_535;

architecture SYN_BEHAVIORAL of FA_535 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_29 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_29;

architecture SYN_rtl of HA_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => A, B => B, Z => S);
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_539 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic);

end FA_539;

architecture SYN_BEHAVIORAL of FA_539 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => A_BAR, B => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_541 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic);

end FA_541;

architecture SYN_BEHAVIORAL of FA_541 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => n6, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => A_BAR, B2 => n1, ZN => Co)
                           ;
   U3 : INV_X1 port map( A => A_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_543 is

   port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic);

end FA_543;

architecture SYN_BEHAVIORAL of FA_543 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n6, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => B_BAR, ZN => Co)
                           ;
   U5 : INV_X1 port map( A => B_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_545 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_545;

architecture SYN_BEHAVIORAL of FA_545 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_546 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_546;

architecture SYN_BEHAVIORAL of FA_546 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1714, n_1715 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG660_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => 
                           n_1714);
   MY_CLK_r_REG654_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1715);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_547 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_547;

architecture SYN_BEHAVIORAL of FA_547 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n7, n8, n9, n11, n12, n_1716 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n4, B => n9, ZN => S);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n9, A2 => n8, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n8, B2 => n9, A => n7, ZN => n3);
   MY_CLK_r_REG664_S1 : DFF_X1 port map( D => A, CK => clk, Q => n9, QN => 
                           n_1716);
   MY_CLK_r_REG666_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n12)
                           ;
   MY_CLK_r_REG356_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n7, QN => n11
                           );
   U1 : XNOR2_X1 port map( A => n11, B => n12, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_548 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_548;

architecture SYN_BEHAVIORAL of FA_548 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n9, n10, n_1717, n_1718 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n9, B => n10, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG667_S1 : DFF_X1 port map( D => B, CK => clk, Q => n10, QN => 
                           n_1717);
   MY_CLK_r_REG342_S1 : DFF_X1 port map( D => n5, CK => clk, Q => n9, QN => 
                           n_1718);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_549 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_549;

architecture SYN_BEHAVIORAL of FA_549 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n6, n7, n_1719, n_1720 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   MY_CLK_r_REG668_S1 : DFF_X1 port map( D => n2, CK => clk, Q => n7, QN => 
                           n_1719);
   MY_CLK_r_REG344_S1 : DFF_X1 port map( D => n3, CK => clk, Q => n6, QN => 
                           n_1720);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_550 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_550;

architecture SYN_BEHAVIORAL of FA_550 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_551 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_551;

architecture SYN_BEHAVIORAL of FA_551 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1721, n_1722 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n8, B => n7, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U3 : XOR2_X1 port map( A => n2, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);
   MY_CLK_r_REG662_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1721);
   MY_CLK_r_REG676_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1722);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_552 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_552;

architecture SYN_BEHAVIORAL of FA_552 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7, n8, n_1723, n_1724 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n7, B => n8, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   MY_CLK_r_REG677_S1 : DFF_X1 port map( D => A, CK => clk, Q => n8, QN => 
                           n_1723);
   MY_CLK_r_REG324_S1 : DFF_X1 port map( D => n4, CK => clk, Q => n7, QN => 
                           n_1724);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_553 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_553;

architecture SYN_BEHAVIORAL of FA_553 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n12, n13, n14, n16, n17, n18 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n8, B => n14, ZN => S);
   U4 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U5 : NAND2_X1 port map( A1 => n14, A2 => n13, ZN => n6);
   U6 : XNOR2_X1 port map( A => n5, B => n4, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n12, A2 => n17, ZN => n5);
   U8 : NAND2_X1 port map( A1 => n12, A2 => n18, ZN => n4);
   MY_CLK_r_REG674_S1 : DFF_X1 port map( D => A, CK => clk, Q => n14, QN => n17
                           );
   MY_CLK_r_REG675_S1 : DFF_X1 port map( D => B, CK => clk, Q => n13, QN => n18
                           );
   MY_CLK_r_REG326_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n12, QN => 
                           n16);
   U1 : XNOR2_X1 port map( A => n16, B => n18, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_554 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_554;

architecture SYN_BEHAVIORAL of FA_554 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n_1725, n_1726 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n7, B => n8, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   MY_CLK_r_REG312_S1 : DFF_X1 port map( D => Ci, CK => clk, Q => n8, QN => 
                           n_1725);
   MY_CLK_r_REG673_S1 : DFF_X1 port map( D => n6, CK => clk, Q => n7, QN => 
                           n_1726);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_555 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_555;

architecture SYN_BEHAVIORAL of FA_555 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28809, net28810, n3, n7, n8, n9, n11, n12, n_1727 : std_logic;

begin
   
   U5 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => net28809);
   U7 : INV_X1 port map( A => Ci, ZN => net28810);
   U2 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   MY_CLK_r_REG316_S1 : DFF_X1 port map( D => net28810, CK => clk, Q => n9, QN 
                           => n_1727);
   MY_CLK_r_REG671_S1 : DFF_X1 port map( D => B, CK => clk, Q => n8, QN => n11)
                           ;
   MY_CLK_r_REG672_S1 : DFF_X1 port map( D => A, CK => clk, Q => n7, QN => n12)
                           ;
   U1 : AOI22_X1 port map( A1 => net28809, A2 => n9, B1 => n12, B2 => n11, ZN 
                           => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_556 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_556;

architecture SYN_BEHAVIORAL of FA_556 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U8 : INV_X1 port map( A => Ci, ZN => n2);
   U2 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n2, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_557 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_557;

architecture SYN_BEHAVIORAL of FA_557 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28819, net28820, net28821, net28822, n5 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => net28821);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net28819);
   U6 : INV_X1 port map( A => B, ZN => net28822);
   U8 : INV_X1 port map( A => Ci, ZN => net28820);
   U9 : AOI22_X1 port map( A1 => net28819, A2 => net28820, B1 => net28821, B2 
                           => net28822, ZN => Co);
   U4 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_558 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_558;

architecture SYN_BEHAVIORAL of FA_558 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U5 : INV_X1 port map( A => A, ZN => n6);
   U6 : INV_X1 port map( A => B, ZN => n5);
   U7 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U8 : INV_X1 port map( A => Ci, ZN => n3);
   U1 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n4, B2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_559 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in std_logic);

end FA_559;

architecture SYN_BEHAVIORAL of FA_559 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net28830, net28833, net28834, n2, n3, n4, n5, n9, n10, n_1728, n_1729
      : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n2, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => Ci, ZN => n2);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net28830);
   U5 : INV_X1 port map( A => B, ZN => net28833);
   U6 : INV_X1 port map( A => A, ZN => net28834);
   U9 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => Co);
   U10 : XNOR2_X1 port map( A => n4, B => n3, ZN => n5);
   U11 : NAND2_X1 port map( A1 => Ci, A2 => net28833, ZN => n3);
   U12 : NAND2_X1 port map( A1 => net28834, A2 => Ci, ZN => n4);
   MY_CLK_r_REG286_S1 : DFF_X1 port map( D => net28830, CK => clk, Q => n10, QN
                           => n_1728);
   MY_CLK_r_REG280_S1 : DFF_X1 port map( D => n5, CK => clk, Q => n9, QN => 
                           n_1729);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_560 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_560;

architecture SYN_BEHAVIORAL of FA_560 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : NOR2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n3);
   U3 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U4 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n2);
   U5 : XNOR2_X1 port map( A => n3, B => A, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_561 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_561;

architecture SYN_BEHAVIORAL of FA_561 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_562 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_562;

architecture SYN_BEHAVIORAL of FA_562 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_563 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_563;

architecture SYN_BEHAVIORAL of FA_563 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_564 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_564;

architecture SYN_BEHAVIORAL of FA_564 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_565 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_565;

architecture SYN_BEHAVIORAL of FA_565 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_566 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_566;

architecture SYN_BEHAVIORAL of FA_566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_568 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_568;

architecture SYN_BEHAVIORAL of FA_568 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n1);
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U6 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_33 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_33;

architecture SYN_rtl of HA_33 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => S);
   U4 : INV_X1 port map( A => A, ZN => n2);
   U5 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);
   U6 : NAND2_X1 port map( A1 => B, A2 => n2, ZN => n3);
   U1 : OR2_X1 port map( A1 => B, A2 => n2, ZN => n4);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_569 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_569;

architecture SYN_BEHAVIORAL of FA_569 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : INV_X1 port map( A => Ci, ZN => n4);
   U5 : INV_X1 port map( A => A, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n2);
   U7 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_570 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_570;

architecture SYN_BEHAVIORAL of FA_570 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U7 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_571 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_571;

architecture SYN_BEHAVIORAL of FA_571 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n8 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U5 : INV_X1 port map( A => A, ZN => n5);
   U6 : INV_X1 port map( A => B, ZN => n4);
   U8 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   U1 : OR2_X1 port map( A1 => A, A2 => B, ZN => n8);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n8, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_572 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_572;

architecture SYN_BEHAVIORAL of FA_572 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_573 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_573;

architecture SYN_BEHAVIORAL of FA_573 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n1);
   U3 : AOI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U6 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_574 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_574;

architecture SYN_BEHAVIORAL of FA_574 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => Ci, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_575 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_575;

architecture SYN_BEHAVIORAL of FA_575 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n5);
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_578 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_578;

architecture SYN_BEHAVIORAL of FA_578 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_579 is

   port( A, B, Ci : in std_logic;  S, Co_BAR : out std_logic);

end FA_579;

architecture SYN_BEHAVIORAL of FA_579 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => Ci, B => n2, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U5 : AND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => Ci, B2 => n3, ZN => Co_BAR
                           );

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_580 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_580;

architecture SYN_BEHAVIORAL of FA_580 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n7, n8 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n2, B => Ci, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n2);
   U5 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U4 : NOR2_X1 port map( A1 => n7, A2 => n3, ZN => Co);
   U6 : NOR2_X1 port map( A1 => Ci, A2 => n8, ZN => n7);
   U7 : AND2_X1 port map( A1 => B, A2 => A, ZN => n8);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_37 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_37;

architecture SYN_rtl of HA_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => B, A2 => n2, ZN => n3);
   U2 : NAND2_X1 port map( A1 => n1, A2 => A, ZN => n4);
   U3 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => S);
   U4 : INV_X1 port map( A => B, ZN => n1);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_38 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_38;

architecture SYN_rtl of HA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_581 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_581;

architecture SYN_BEHAVIORAL of FA_581 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n3, A2 => n4, B1 => n2, B2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_582 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_582;

architecture SYN_BEHAVIORAL of FA_582 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => B, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_583 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_583;

architecture SYN_BEHAVIORAL of FA_583 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4 : std_logic;

begin
   
   U2 : NAND2_X1 port map( A1 => n3, A2 => n2, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => n4, ZN => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n2);
   U5 : XNOR2_X1 port map( A => Ci, B => B, ZN => n4);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_584 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_584;

architecture SYN_BEHAVIORAL of FA_584 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U2 : INV_X1 port map( A => A, ZN => n2);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_585 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_585;

architecture SYN_BEHAVIORAL of FA_585 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_586 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_586;

architecture SYN_BEHAVIORAL of FA_586 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n8 : std_logic;

begin
   
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => A, ZN => n2);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U2 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U7 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U8 : XNOR2_X1 port map( A => n8, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_587 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_587;

architecture SYN_BEHAVIORAL of FA_587 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n7 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n4);
   U5 : INV_X1 port map( A => B, ZN => n3);
   U6 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);
   U7 : OAI21_X1 port map( B1 => n4, B2 => n3, A => n2, ZN => Co);
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U2 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_588 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_588;

architecture SYN_BEHAVIORAL of FA_588 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_589 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_589;

architecture SYN_BEHAVIORAL of FA_589 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U2 : XNOR2_X1 port map( A => n5, B => A, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => A, ZN => n2);
   U7 : INV_X1 port map( A => B, ZN => n1);
   U1 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n1, B2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_590 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_590;

architecture SYN_BEHAVIORAL of FA_590 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n6 : std_logic;

begin
   
   U2 : INV_X1 port map( A => Ci, ZN => n2);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U4 : NOR2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U5 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U1 : AOI21_X1 port map( B1 => n2, B2 => n3, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_591 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_591;

architecture SYN_BEHAVIORAL of FA_591 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n1, B => A, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => B, ZN => n1);
   U3 : NOR2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U5 : AOI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n6);
   U4 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_592 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_592;

architecture SYN_BEHAVIORAL of FA_592 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n1, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => Ci, ZN => n1);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);
   U5 : OAI21_X1 port map( B1 => A, B2 => B, A => Ci, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_40 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_40;

architecture SYN_rtl of HA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_41 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_41;

architecture SYN_rtl of HA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_42 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_42;

architecture SYN_rtl of HA_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   C <= B;
   
   U1 : INV_X1 port map( A => B, ZN => S);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_593 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_593;

architecture SYN_BEHAVIORAL of FA_593 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_594 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_594;

architecture SYN_BEHAVIORAL of FA_594 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_595 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_595;

architecture SYN_BEHAVIORAL of FA_595 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n1);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n2);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_596 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_596;

architecture SYN_BEHAVIORAL of FA_596 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U5 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U1 : OAI21_X1 port map( B1 => B, B2 => n3, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_597 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic);

end FA_597;

architecture SYN_BEHAVIORAL of FA_597 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n5, ZN => S);
   U2 : XNOR2_X1 port map( A => n7, B => Ci, ZN => n5);
   U3 : NAND2_X1 port map( A1 => B, A2 => n7, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : INV_X1 port map( A => B, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => A_BAR, B2 => n1, ZN => Co)
                           ;
   U5 : INV_X1 port map( A => A_BAR, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_598 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_598;

architecture SYN_BEHAVIORAL of FA_598 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U2 : INV_X1 port map( A => B, ZN => n2);
   U1 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => Co);
   U3 : XNOR2_X1 port map( A => Ci, B => B, ZN => S);
   U4 : INV_X1 port map( A => Ci, ZN => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_599 is

   port( Ci : in std_logic;  S, Co : out std_logic;  B_BAR, A_BAR : in 
         std_logic);

end FA_599;

architecture SYN_BEHAVIORAL of FA_599 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => A_BAR, B => n6, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => A_BAR, B2 => B_BAR, ZN => 
                           Co);
   U5 : INV_X1 port map( A => B_BAR, ZN => n6);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_600 is

   port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic);

end FA_600;

architecture SYN_BEHAVIORAL of FA_600 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XOR2_X1 port map( A => A_BAR, B => B, Z => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n3);
   U5 : INV_X1 port map( A => B, ZN => n1);
   U6 : OAI22_X1 port map( A1 => n4, A2 => n3, B1 => A_BAR, B2 => n1, ZN => Co)
                           ;

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_601 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_601;

architecture SYN_BEHAVIORAL of FA_601 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n4, ZN => S);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n4);
   U3 : INV_X1 port map( A => A, ZN => n3);
   U4 : INV_X1 port map( A => B, ZN => n2);
   U5 : OAI21_X1 port map( B1 => B, B2 => A, A => Ci, ZN => n1);
   U6 : OAI21_X1 port map( B1 => n3, B2 => n2, A => n1, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_602 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_602;

architecture SYN_BEHAVIORAL of FA_602 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n1);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n2);
   U4 : XNOR2_X1 port map( A => B, B => n7, ZN => S);
   U5 : XNOR2_X1 port map( A => Ci, B => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U7 : INV_X1 port map( A => Ci, ZN => n5);
   U8 : INV_X1 port map( A => A, ZN => n4);
   U9 : INV_X1 port map( A => B, ZN => n3);
   U3 : AND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_603 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_603;

architecture SYN_BEHAVIORAL of FA_603 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29038, net29039, net29040, n1, n2, n3, n4 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);
   U3 : NAND2_X1 port map( A1 => n4, A2 => net29038, ZN => n1);
   U4 : NAND2_X1 port map( A1 => net29039, A2 => net29040, ZN => n2);
   U5 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U7 : INV_X1 port map( A => Ci, ZN => net29038);
   U8 : INV_X1 port map( A => A, ZN => net29039);
   U9 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U10 : INV_X1 port map( A => B, ZN => net29040);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_604 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_604;

architecture SYN_BEHAVIORAL of FA_604 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n7 : std_logic;

begin
   
   U3 : INV_X1 port map( A => A, ZN => n4);
   U4 : INV_X1 port map( A => B, ZN => n3);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n2);
   U6 : INV_X1 port map( A => Ci, ZN => n1);
   U7 : AOI22_X1 port map( A1 => n4, A2 => n3, B1 => n2, B2 => n1, ZN => Co);
   U2 : XNOR2_X1 port map( A => Ci, B => A, ZN => n7);
   U1 : XNOR2_X1 port map( A => n7, B => B, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_605 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_605;

architecture SYN_BEHAVIORAL of FA_605 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U2 : INV_X1 port map( A => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => n2);
   U7 : XNOR2_X1 port map( A => n9, B => Ci, ZN => S);
   U8 : XNOR2_X1 port map( A => B, B => A, ZN => n9);
   U9 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n8);
   U10 : INV_X1 port map( A => Ci, ZN => n7);
   U11 : INV_X1 port map( A => B, ZN => n5);
   U5 : AND2_X1 port map( A1 => n1, A2 => n2, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_606 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_606;

architecture SYN_BEHAVIORAL of FA_606 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n9 : std_logic;

begin
   
   U5 : INV_X1 port map( A => A, ZN => n6);
   U6 : INV_X1 port map( A => B, ZN => n5);
   U7 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U8 : INV_X1 port map( A => Ci, ZN => n3);
   U1 : AOI22_X1 port map( A1 => n6, A2 => n5, B1 => n3, B2 => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => Ci, B => n9, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n9);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_607 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_607;

architecture SYN_BEHAVIORAL of FA_607 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29057, net29058, n7, n8, n9, n10 : std_logic;

begin
   
   U8 : INV_X1 port map( A => A, ZN => net29057);
   U10 : INV_X1 port map( A => B, ZN => net29058);
   U1 : NOR2_X1 port map( A1 => n7, A2 => Ci, ZN => n8);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => n7);
   U3 : NOR2_X1 port map( A1 => n8, A2 => n9, ZN => Co);
   U4 : AND2_X1 port map( A1 => net29057, A2 => net29058, ZN => n9);
   U5 : XNOR2_X1 port map( A => Ci, B => n10, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n10);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n7 : std_logic;

begin
   
   U4 : INV_X1 port map( A => A, ZN => n5);
   U5 : INV_X1 port map( A => B, ZN => n4);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n3);
   U7 : INV_X1 port map( A => Ci, ZN => n2);
   U1 : AOI22_X1 port map( A1 => n5, A2 => n4, B1 => n3, B2 => n2, ZN => Co);
   U2 : XNOR2_X1 port map( A => n7, B => B, ZN => S);
   U3 : XNOR2_X1 port map( A => Ci, B => A, ZN => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_43 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_43;

architecture SYN_rtl of HA_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => B, B => A, Z => S);
   U1 : AND2_X1 port map( A1 => A, A2 => B, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity HA_0 is

   port( A, B : in std_logic;  S, C : out std_logic);

end HA_0;

architecture SYN_rtl of HA_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => A, B => B, Z => S);
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => C);

end SYN_rtl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_5 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
         p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
         p_23_port, p_18_BAR, p_12_port, p_11_port, p_10_port, p_9_port, 
         p_8_port, p_6_port, p_3_port, p_1_port, p_0_port, p_17_BAR, p_20_BAR, 
         p_19_BAR, p_22_BAR, p_21_BAR, p_7_BAR, p_5_BAR, p_4_BAR, p_2_BAR, 
         p_14_BAR, p_13_BAR, p_16_BAR, p_15_BAR : out std_logic);

end ENC_5;

architecture SYN_beh of ENC_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U3 : NAND2_X1 port map( A1 => A(7), A2 => b(0), ZN => p_7_BAR);
   U4 : NAND2_X1 port map( A1 => A(2), A2 => b(0), ZN => p_2_BAR);
   U5 : NAND2_X1 port map( A1 => A(20), A2 => b(0), ZN => p_20_BAR);
   U6 : NAND2_X1 port map( A1 => A(4), A2 => b(0), ZN => p_4_BAR);
   U7 : NAND2_X1 port map( A1 => A(5), A2 => b(0), ZN => p_5_BAR);
   U9 : AND2_X1 port map( A1 => A(12), A2 => b(0), ZN => p_12_port);
   U10 : AND2_X1 port map( A1 => A(11), A2 => b(0), ZN => p_11_port);
   U11 : AND2_X1 port map( A1 => A(1), A2 => b(0), ZN => p_1_port);
   U12 : AND2_X1 port map( A1 => A(0), A2 => b(0), ZN => p_0_port);
   U13 : AND2_X1 port map( A1 => A(23), A2 => b(0), ZN => p_23_port);
   U14 : AND2_X1 port map( A1 => A(6), A2 => b(0), ZN => p_6_port);
   U15 : AND2_X1 port map( A1 => A(3), A2 => b(0), ZN => p_3_port);
   U16 : AND2_X1 port map( A1 => A(10), A2 => b(0), ZN => p_10_port);
   U17 : AND2_X1 port map( A1 => A(9), A2 => b(0), ZN => p_9_port);
   U18 : AND2_X1 port map( A1 => A(8), A2 => b(0), ZN => p_8_port);
   U20 : NAND2_X1 port map( A1 => A(22), A2 => b(0), ZN => p_22_BAR);
   U21 : NAND2_X1 port map( A1 => A(21), A2 => b(0), ZN => p_21_BAR);
   U22 : NAND2_X1 port map( A1 => A(19), A2 => b(0), ZN => p_19_BAR);
   U23 : NAND2_X1 port map( A1 => A(18), A2 => b(0), ZN => p_18_BAR);
   U24 : NAND2_X1 port map( A1 => A(17), A2 => b(0), ZN => p_17_BAR);
   U25 : NAND2_X1 port map( A1 => A(16), A2 => b(0), ZN => p_16_BAR);
   U26 : NAND2_X1 port map( A1 => A(15), A2 => b(0), ZN => p_15_BAR);
   U27 : NAND2_X1 port map( A1 => A(14), A2 => b(0), ZN => p_14_BAR);
   U29 : NAND2_X1 port map( A1 => A(13), A2 => b(0), ZN => p_13_BAR);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_6 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_6;

architecture SYN_beh of ENC_6 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29488, net29492, net29502, net29521, net29523, net31045, net29525,
      net29490, net29455, net29452, net29451, n3, n4, n5, n6, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n56, n60
      , n63, n64, n65, n66, n71, n72 : std_logic;

begin
   
   U9 : NAND3_X1 port map( A1 => n5, A2 => net29455, A3 => net29490, ZN => 
                           p(14));
   U10 : MUX2_X1 port map( A => n72, B => net29451, S => A(14), Z => net29488);
   U11 : MUX2_X1 port map( A => n65, B => net31045, S => A(14), Z => n5);
   U12 : XNOR2_X1 port map( A => b(1), B => b(0), ZN => n4);
   U13 : OR2_X1 port map( A1 => b(1), A2 => b(0), ZN => n6);
   U18 : MUX2_X1 port map( A => n64, B => net29451, S => A(13), Z => net29490);
   U23 : MUX2_X1 port map( A => n66, B => net31045, S => A(13), Z => net29492);
   U29 : INV_X1 port map( A => b(0), ZN => net29525);
   U30 : MUX2_X1 port map( A => net29521, B => net31045, S => A(0), Z => 
                           net29523);
   U39 : INV_X1 port map( A => b(2), ZN => net29502);
   U41 : NAND2_X1 port map( A1 => b(2), A2 => n10, ZN => net29521);
   U42 : OAI211_X1 port map( C1 => net29502, C2 => n10, A => net29452, B => 
                           net29523, ZN => p(0));
   U43 : MUX2_X1 port map( A => n72, B => net29451, S => A(0), Z => n12);
   U44 : MUX2_X1 port map( A => n66, B => net31045, S => A(1), Z => n11);
   U45 : NAND3_X1 port map( A1 => n12, A2 => n63, A3 => n11, ZN => p(1));
   U46 : MUX2_X1 port map( A => n64, B => net29451, S => A(1), Z => n14);
   U47 : MUX2_X1 port map( A => n65, B => net31045, S => A(2), Z => n13);
   U48 : NAND3_X1 port map( A1 => n13, A2 => n63, A3 => n14, ZN => p(2));
   U49 : MUX2_X1 port map( A => n71, B => net29451, S => A(2), Z => n16);
   U50 : MUX2_X1 port map( A => n65, B => net31045, S => A(3), Z => n15);
   U51 : NAND3_X1 port map( A1 => n16, A2 => net29455, A3 => n15, ZN => p(3));
   U52 : MUX2_X1 port map( A => n64, B => net29451, S => A(3), Z => n18);
   U53 : MUX2_X1 port map( A => n66, B => net31045, S => A(4), Z => n17);
   U54 : NAND3_X1 port map( A1 => n17, A2 => n63, A3 => n18, ZN => p(4));
   U55 : MUX2_X1 port map( A => n66, B => net31045, S => A(5), Z => n20);
   U56 : MUX2_X1 port map( A => n64, B => net29451, S => A(4), Z => n19);
   U57 : NAND3_X1 port map( A1 => n20, A2 => n63, A3 => n19, ZN => p(5));
   U58 : MUX2_X1 port map( A => n71, B => net29451, S => A(5), Z => n22);
   U59 : MUX2_X1 port map( A => n65, B => net31045, S => A(6), Z => n21);
   U60 : NAND3_X1 port map( A1 => n22, A2 => n63, A3 => n21, ZN => p(6));
   U61 : MUX2_X1 port map( A => n72, B => net29451, S => A(6), Z => n24);
   U62 : MUX2_X1 port map( A => n66, B => net31045, S => A(7), Z => n23);
   U63 : NAND3_X1 port map( A1 => n24, A2 => n63, A3 => n23, ZN => p(7));
   U64 : MUX2_X1 port map( A => n72, B => net29451, S => A(7), Z => n26);
   U65 : MUX2_X1 port map( A => n66, B => net31045, S => A(8), Z => n25);
   U66 : NAND3_X1 port map( A1 => n26, A2 => n25, A3 => net29455, ZN => p(8));
   U67 : MUX2_X1 port map( A => n72, B => net29451, S => A(8), Z => n28);
   U68 : MUX2_X1 port map( A => n65, B => net31045, S => A(9), Z => n27);
   U69 : NAND3_X1 port map( A1 => n28, A2 => net29455, A3 => n27, ZN => p(9));
   U70 : MUX2_X1 port map( A => n64, B => net29451, S => A(9), Z => n32);
   U71 : XOR2_X1 port map( A => b(1), B => b(0), Z => n29);
   U72 : NAND2_X1 port map( A1 => n29, A2 => net29502, ZN => n30);
   U73 : MUX2_X1 port map( A => n66, B => n30, S => A(10), Z => n31);
   U74 : NAND3_X1 port map( A1 => net29455, A2 => n32, A3 => n31, ZN => p(10));
   U75 : MUX2_X1 port map( A => net29452, B => net29451, S => A(10), Z => n34);
   U76 : MUX2_X1 port map( A => n66, B => net31045, S => A(11), Z => n33);
   U77 : NAND3_X1 port map( A1 => n34, A2 => net29455, A3 => n33, ZN => p(11));
   U78 : MUX2_X1 port map( A => n64, B => net29451, S => A(11), Z => n36);
   U79 : MUX2_X1 port map( A => n66, B => net31045, S => A(12), Z => n35);
   U80 : NAND3_X1 port map( A1 => n36, A2 => net29455, A3 => n35, ZN => p(12));
   U81 : MUX2_X1 port map( A => n64, B => net29451, S => A(12), Z => n37);
   U82 : NAND3_X1 port map( A1 => net29492, A2 => n37, A3 => net29455, ZN => 
                           p(13));
   U83 : MUX2_X1 port map( A => n66, B => net31045, S => A(15), Z => n38);
   U84 : NAND3_X1 port map( A1 => net29488, A2 => net29455, A3 => n38, ZN => 
                           p(15));
   U85 : MUX2_X1 port map( A => n64, B => net29451, S => A(15), Z => n40);
   U86 : MUX2_X1 port map( A => n66, B => net31045, S => A(16), Z => n39);
   U87 : NAND3_X1 port map( A1 => n40, A2 => net29455, A3 => n39, ZN => p(16));
   U88 : MUX2_X1 port map( A => n71, B => net29451, S => A(16), Z => n42);
   U89 : MUX2_X1 port map( A => n65, B => net31045, S => A(17), Z => n41);
   U90 : NAND3_X1 port map( A1 => n42, A2 => net29455, A3 => n41, ZN => p(17));
   U91 : MUX2_X1 port map( A => net29452, B => net29451, S => A(17), Z => n44);
   U92 : MUX2_X1 port map( A => n65, B => net31045, S => A(18), Z => n43);
   U93 : NAND3_X1 port map( A1 => n44, A2 => net29455, A3 => n43, ZN => p(18));
   U94 : MUX2_X1 port map( A => n66, B => net31045, S => A(19), Z => n46);
   U95 : MUX2_X1 port map( A => n64, B => net29451, S => A(18), Z => n45);
   U96 : NAND3_X1 port map( A1 => n63, A2 => n46, A3 => n45, ZN => p(19));
   U97 : MUX2_X1 port map( A => net29452, B => net29451, S => A(19), Z => n48);
   U98 : MUX2_X1 port map( A => n65, B => net31045, S => A(20), Z => n47);
   U99 : NAND3_X1 port map( A1 => n48, A2 => n63, A3 => n47, ZN => p(20));
   U100 : MUX2_X1 port map( A => n71, B => net29451, S => A(20), Z => n50);
   U101 : MUX2_X1 port map( A => n65, B => net31045, S => A(21), Z => n49);
   U102 : NAND3_X1 port map( A1 => n50, A2 => net29455, A3 => n49, ZN => p(21))
                           ;
   U103 : MUX2_X1 port map( A => n71, B => net29451, S => A(21), Z => n52);
   U104 : MUX2_X1 port map( A => n65, B => net31045, S => A(22), Z => n51);
   U105 : NAND3_X1 port map( A1 => n52, A2 => n63, A3 => n51, ZN => p(22));
   U106 : MUX2_X1 port map( A => n64, B => n10, S => A(22), Z => n54);
   U107 : MUX2_X1 port map( A => n65, B => net31045, S => A(23), Z => n53);
   U108 : NAND3_X1 port map( A1 => n54, A2 => n63, A3 => n53, ZN => p(23));
   U109 : MUX2_X1 port map( A => n71, B => net29451, S => A(23), Z => n56);
   U111 : NAND3_X1 port map( A1 => n56, A2 => n63, A3 => n65, ZN => p(24));
   U114 : NAND3_X1 port map( A1 => net29452, A2 => n63, A3 => n65, ZN => p(25))
                           ;
   U8 : OR2_X2 port map( A1 => b(2), A2 => n4, ZN => net31045);
   U16 : NAND3_X1 port map( A1 => b(2), A2 => net29525, A3 => n60, ZN => n64);
   U20 : NAND2_X1 port map( A1 => n6, A2 => b(2), ZN => n3);
   U4 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => net29451);
   U3 : NAND2_X2 port map( A1 => b(2), A2 => net29521, ZN => net29455);
   U6 : NAND2_X2 port map( A1 => b(2), A2 => net29521, ZN => n63);
   U7 : CLKBUF_X2 port map( A => n3, Z => n66);
   U14 : CLKBUF_X2 port map( A => n3, Z => n65);
   U15 : INV_X1 port map( A => b(1), ZN => n60);
   U17 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n10);
   U19 : NAND3_X1 port map( A1 => b(2), A2 => net29525, A3 => n60, ZN => n71);
   U21 : NAND3_X1 port map( A1 => b(2), A2 => net29525, A3 => n60, ZN => n72);
   U22 : NAND3_X1 port map( A1 => b(2), A2 => net29525, A3 => n60, ZN => 
                           net29452);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_7 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_7;

architecture SYN_beh of ENC_7 is

   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n85, n87, n89, n90
      , n91, n18, n71 : std_logic;

begin
   
   U3 : NAND3_X1 port map( A1 => n56, A2 => n87, A3 => n55, ZN => p(16));
   U4 : OR2_X1 port map( A1 => n20, A2 => b(2), ZN => n1);
   U24 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n20);
   U27 : INV_X1 port map( A => b(2), ZN => n23);
   U28 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n22);
   U29 : INV_X1 port map( A => b(0), ZN => n19);
   U32 : NAND2_X1 port map( A1 => b(2), A2 => n22, ZN => n24);
   U33 : MUX2_X1 port map( A => n24, B => n1, S => A(0), Z => n21);
   U34 : OAI211_X1 port map( C1 => n23, C2 => n22, A => n90, B => n21, ZN => 
                           p(0));
   U36 : MUX2_X1 port map( A => n90, B => n91, S => A(0), Z => n26);
   U39 : MUX2_X1 port map( A => n89, B => n85, S => A(1), Z => n25);
   U40 : NAND3_X1 port map( A1 => n26, A2 => n87, A3 => n25, ZN => p(1));
   U41 : MUX2_X1 port map( A => n90, B => n91, S => A(1), Z => n28);
   U42 : MUX2_X1 port map( A => n89, B => n85, S => A(2), Z => n27);
   U43 : NAND3_X1 port map( A1 => n28, A2 => n87, A3 => n27, ZN => p(2));
   U44 : MUX2_X1 port map( A => n90, B => n91, S => A(2), Z => n30);
   U45 : MUX2_X1 port map( A => n89, B => n85, S => A(3), Z => n29);
   U46 : NAND3_X1 port map( A1 => n30, A2 => n87, A3 => n29, ZN => p(3));
   U47 : MUX2_X1 port map( A => n90, B => n91, S => A(3), Z => n32);
   U48 : MUX2_X1 port map( A => n89, B => n85, S => A(4), Z => n31);
   U49 : NAND3_X1 port map( A1 => n32, A2 => n87, A3 => n31, ZN => p(4));
   U50 : MUX2_X1 port map( A => n89, B => n85, S => A(5), Z => n34);
   U51 : MUX2_X1 port map( A => n90, B => n91, S => A(4), Z => n33);
   U52 : NAND3_X1 port map( A1 => n34, A2 => n87, A3 => n33, ZN => p(5));
   U53 : MUX2_X1 port map( A => n90, B => n91, S => A(5), Z => n36);
   U54 : MUX2_X1 port map( A => n89, B => n1, S => A(6), Z => n35);
   U55 : NAND3_X1 port map( A1 => n36, A2 => n87, A3 => n35, ZN => p(6));
   U56 : MUX2_X1 port map( A => n90, B => n91, S => A(6), Z => n38);
   U57 : MUX2_X1 port map( A => n89, B => n85, S => A(7), Z => n37);
   U58 : NAND3_X1 port map( A1 => n38, A2 => n87, A3 => n37, ZN => p(7));
   U59 : MUX2_X1 port map( A => n89, B => n85, S => A(8), Z => n40);
   U60 : MUX2_X1 port map( A => n90, B => n91, S => A(7), Z => n39);
   U61 : NAND3_X1 port map( A1 => n87, A2 => n40, A3 => n39, ZN => p(8));
   U62 : MUX2_X1 port map( A => n90, B => n91, S => A(8), Z => n42);
   U63 : MUX2_X1 port map( A => n89, B => n1, S => A(9), Z => n41);
   U64 : NAND3_X1 port map( A1 => n42, A2 => n87, A3 => n41, ZN => p(9));
   U65 : MUX2_X1 port map( A => n90, B => n91, S => A(9), Z => n44);
   U66 : MUX2_X1 port map( A => n89, B => n85, S => A(10), Z => n43);
   U67 : NAND3_X1 port map( A1 => n44, A2 => n87, A3 => n43, ZN => p(10));
   U68 : MUX2_X1 port map( A => n89, B => n1, S => A(11), Z => n46);
   U69 : MUX2_X1 port map( A => n90, B => n91, S => A(10), Z => n45);
   U70 : NAND3_X1 port map( A1 => n46, A2 => n45, A3 => n87, ZN => p(11));
   U71 : MUX2_X1 port map( A => n89, B => n1, S => A(12), Z => n48);
   U72 : MUX2_X1 port map( A => n90, B => n91, S => A(11), Z => n47);
   U73 : NAND3_X1 port map( A1 => n48, A2 => n47, A3 => n87, ZN => p(12));
   U74 : MUX2_X1 port map( A => n90, B => n91, S => A(12), Z => n50);
   U75 : MUX2_X1 port map( A => n89, B => n1, S => A(13), Z => n49);
   U76 : NAND3_X1 port map( A1 => n50, A2 => n87, A3 => n49, ZN => p(13));
   U77 : MUX2_X1 port map( A => n90, B => n91, S => A(13), Z => n52);
   U78 : MUX2_X1 port map( A => n89, B => n85, S => A(14), Z => n51);
   U79 : NAND3_X1 port map( A1 => n52, A2 => n87, A3 => n51, ZN => p(14));
   U80 : MUX2_X1 port map( A => n90, B => n91, S => A(14), Z => n54);
   U81 : MUX2_X1 port map( A => n89, B => n1, S => A(15), Z => n53);
   U82 : NAND3_X1 port map( A1 => n54, A2 => n87, A3 => n53, ZN => p(15));
   U83 : MUX2_X1 port map( A => n90, B => n91, S => A(15), Z => n56);
   U84 : MUX2_X1 port map( A => n89, B => n85, S => A(16), Z => n55);
   U85 : MUX2_X1 port map( A => n90, B => n91, S => A(16), Z => n58);
   U86 : MUX2_X1 port map( A => n89, B => n85, S => A(17), Z => n57);
   U87 : NAND3_X1 port map( A1 => n58, A2 => n87, A3 => n57, ZN => p(17));
   U88 : MUX2_X1 port map( A => n90, B => n91, S => A(17), Z => n60);
   U89 : MUX2_X1 port map( A => n89, B => n85, S => A(18), Z => n59);
   U90 : NAND3_X1 port map( A1 => n60, A2 => n87, A3 => n59, ZN => p(18));
   U91 : MUX2_X1 port map( A => n90, B => n91, S => A(18), Z => n62);
   U92 : MUX2_X1 port map( A => n89, B => n85, S => A(19), Z => n61);
   U93 : NAND3_X1 port map( A1 => n62, A2 => n87, A3 => n61, ZN => p(19));
   U94 : MUX2_X1 port map( A => n90, B => n91, S => A(19), Z => n64);
   U95 : MUX2_X1 port map( A => n89, B => n1, S => A(20), Z => n63);
   U96 : NAND3_X1 port map( A1 => n64, A2 => n87, A3 => n63, ZN => p(20));
   U97 : MUX2_X1 port map( A => n90, B => n91, S => A(20), Z => n66);
   U98 : MUX2_X1 port map( A => n89, B => n85, S => A(21), Z => n65);
   U99 : NAND3_X1 port map( A1 => n66, A2 => n87, A3 => n65, ZN => p(21));
   U100 : MUX2_X1 port map( A => n90, B => n91, S => A(21), Z => n68);
   U101 : MUX2_X1 port map( A => n89, B => n85, S => A(22), Z => n67);
   U102 : NAND3_X1 port map( A1 => n68, A2 => n87, A3 => n67, ZN => p(22));
   U103 : MUX2_X1 port map( A => n90, B => n91, S => A(22), Z => n70);
   U104 : MUX2_X1 port map( A => n89, B => n85, S => A(23), Z => n69);
   U105 : NAND3_X1 port map( A1 => n70, A2 => n87, A3 => n69, ZN => p(23));
   U106 : MUX2_X1 port map( A => n90, B => n91, S => A(23), Z => n72);
   U108 : NAND3_X1 port map( A1 => n72, A2 => n87, A3 => n89, ZN => p(24));
   U114 : NAND3_X1 port map( A1 => n90, A2 => n87, A3 => n89, ZN => p(26));
   U117 : NAND3_X1 port map( A1 => n90, A2 => n87, A3 => n89, ZN => p(27));
   U6 : OR2_X1 port map( A1 => n20, A2 => b(2), ZN => n85);
   U11 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n91);
   U111 : NAND3_X1 port map( A1 => n90, A2 => n87, A3 => n89, ZN => p(25));
   U37 : NAND2_X2 port map( A1 => b(2), A2 => n24, ZN => n87);
   U5 : NAND2_X2 port map( A1 => b(2), A2 => n71, ZN => n89);
   U7 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n71);
   U8 : INV_X1 port map( A => b(1), ZN => n18);
   U9 : NAND3_X2 port map( A1 => b(2), A2 => n19, A3 => n18, ZN => n90);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_8 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_8;

architecture SYN_beh of ENC_8 is

   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal p_29_port, p_28_port, p_26_port, p_25_port, p_24_port, p_23_port, 
      p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, p_17_port, 
      p_16_port, p_15_port, p_14_port, p_13_port, p_12_port, p_11_port, 
      p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, p_5_port, p_4_port, 
      p_3_port, p_2_port, p_1_port, p_0_port, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, 
      n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54
      , n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, 
      n69, n71, n84, n86, n88, n89, n90, n17, n73, n77, n78, n_1789, n_1790, 
      n_1791 : std_logic;

begin
   p <= ( n_1789, n_1790, n_1791, p_29_port, p_28_port, p_28_port, p_26_port, 
      p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, p_20_port, 
      p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, p_14_port, 
      p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port, p_7_port,
      p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, p_0_port );
   
   U20 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n19);
   U23 : INV_X1 port map( A => b(2), ZN => n22);
   U24 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n21);
   U28 : NAND2_X1 port map( A1 => b(2), A2 => n21, ZN => n23);
   U29 : MUX2_X1 port map( A => n23, B => n84, S => A(0), Z => n20);
   U30 : OAI211_X1 port map( C1 => n22, C2 => n21, A => n77, B => n20, ZN => 
                           p_0_port);
   U32 : MUX2_X1 port map( A => n78, B => n90, S => A(0), Z => n25);
   U35 : MUX2_X1 port map( A => n88, B => n84, S => A(1), Z => n24);
   U36 : NAND3_X1 port map( A1 => n25, A2 => n86, A3 => n24, ZN => p_1_port);
   U37 : MUX2_X1 port map( A => n78, B => n90, S => A(1), Z => n27);
   U38 : MUX2_X1 port map( A => n88, B => n84, S => A(2), Z => n26);
   U39 : NAND3_X1 port map( A1 => n27, A2 => n86, A3 => n26, ZN => p_2_port);
   U40 : MUX2_X1 port map( A => n78, B => n90, S => A(2), Z => n29);
   U41 : MUX2_X1 port map( A => n88, B => n84, S => A(3), Z => n28);
   U42 : NAND3_X1 port map( A1 => n29, A2 => n86, A3 => n28, ZN => p_3_port);
   U43 : MUX2_X1 port map( A => n77, B => n90, S => A(3), Z => n31);
   U44 : MUX2_X1 port map( A => n88, B => n84, S => A(4), Z => n30);
   U45 : NAND3_X1 port map( A1 => n31, A2 => n86, A3 => n30, ZN => p_4_port);
   U46 : MUX2_X1 port map( A => n77, B => n90, S => A(4), Z => n33);
   U47 : MUX2_X1 port map( A => n88, B => n84, S => A(5), Z => n32);
   U48 : NAND3_X1 port map( A1 => n33, A2 => n86, A3 => n32, ZN => p_5_port);
   U49 : MUX2_X1 port map( A => n78, B => n90, S => A(5), Z => n35);
   U50 : MUX2_X1 port map( A => n88, B => n84, S => A(6), Z => n34);
   U51 : NAND3_X1 port map( A1 => n35, A2 => n86, A3 => n34, ZN => p_6_port);
   U52 : MUX2_X1 port map( A => n88, B => n84, S => A(7), Z => n37);
   U53 : MUX2_X1 port map( A => n78, B => n90, S => A(6), Z => n36);
   U54 : NAND3_X1 port map( A1 => n37, A2 => n86, A3 => n36, ZN => p_7_port);
   U55 : MUX2_X1 port map( A => n88, B => n84, S => A(8), Z => n39);
   U56 : MUX2_X1 port map( A => n78, B => n90, S => A(7), Z => n38);
   U57 : NAND3_X1 port map( A1 => n39, A2 => n86, A3 => n38, ZN => p_8_port);
   U58 : MUX2_X1 port map( A => n77, B => n90, S => A(8), Z => n41);
   U59 : MUX2_X1 port map( A => n88, B => n84, S => A(9), Z => n40);
   U60 : NAND3_X1 port map( A1 => n41, A2 => n86, A3 => n40, ZN => p_9_port);
   U61 : MUX2_X1 port map( A => n88, B => n84, S => A(10), Z => n43);
   U62 : MUX2_X1 port map( A => n77, B => n90, S => A(9), Z => n42);
   U63 : NAND3_X1 port map( A1 => n86, A2 => n43, A3 => n42, ZN => p_10_port);
   U64 : MUX2_X1 port map( A => n77, B => n90, S => A(10), Z => n45);
   U65 : MUX2_X1 port map( A => n88, B => n84, S => A(11), Z => n44);
   U66 : NAND3_X1 port map( A1 => n45, A2 => n86, A3 => n44, ZN => p_11_port);
   U67 : MUX2_X1 port map( A => n78, B => n90, S => A(11), Z => n47);
   U68 : MUX2_X1 port map( A => n88, B => n84, S => A(12), Z => n46);
   U69 : NAND3_X1 port map( A1 => n47, A2 => n86, A3 => n46, ZN => p_12_port);
   U70 : MUX2_X1 port map( A => n88, B => n84, S => A(13), Z => n49);
   U71 : MUX2_X1 port map( A => n77, B => n90, S => A(12), Z => n48);
   U72 : NAND3_X1 port map( A1 => n49, A2 => n86, A3 => n48, ZN => p_13_port);
   U73 : MUX2_X1 port map( A => n88, B => n84, S => A(14), Z => n51);
   U74 : MUX2_X1 port map( A => n77, B => n90, S => A(13), Z => n50);
   U75 : NAND3_X1 port map( A1 => n51, A2 => n50, A3 => n86, ZN => p_14_port);
   U76 : MUX2_X1 port map( A => n77, B => n90, S => A(14), Z => n53);
   U77 : MUX2_X1 port map( A => n88, B => n84, S => A(15), Z => n52);
   U78 : NAND3_X1 port map( A1 => n52, A2 => n53, A3 => n86, ZN => p_15_port);
   U79 : MUX2_X1 port map( A => n88, B => n84, S => A(16), Z => n55);
   U80 : MUX2_X1 port map( A => n89, B => n90, S => A(15), Z => n54);
   U81 : NAND3_X1 port map( A1 => n55, A2 => n86, A3 => n54, ZN => p_16_port);
   U82 : MUX2_X1 port map( A => n77, B => n90, S => A(16), Z => n57);
   U83 : MUX2_X1 port map( A => n88, B => n84, S => A(17), Z => n56);
   U84 : NAND3_X1 port map( A1 => n57, A2 => n86, A3 => n56, ZN => p_17_port);
   U85 : MUX2_X1 port map( A => n77, B => n90, S => A(17), Z => n59);
   U86 : MUX2_X1 port map( A => n88, B => n84, S => A(18), Z => n58);
   U87 : NAND3_X1 port map( A1 => n58, A2 => n86, A3 => n59, ZN => p_18_port);
   U88 : MUX2_X1 port map( A => n78, B => n90, S => A(18), Z => n61);
   U89 : MUX2_X1 port map( A => n88, B => n84, S => A(19), Z => n60);
   U90 : NAND3_X1 port map( A1 => n61, A2 => n86, A3 => n60, ZN => p_19_port);
   U91 : MUX2_X1 port map( A => n77, B => n90, S => A(19), Z => n63);
   U92 : MUX2_X1 port map( A => n88, B => n84, S => A(20), Z => n62);
   U93 : NAND3_X1 port map( A1 => n63, A2 => n86, A3 => n62, ZN => p_20_port);
   U94 : MUX2_X1 port map( A => n78, B => n90, S => A(20), Z => n65);
   U95 : MUX2_X1 port map( A => n88, B => n84, S => A(21), Z => n64);
   U96 : NAND3_X1 port map( A1 => n65, A2 => n86, A3 => n64, ZN => p_21_port);
   U97 : MUX2_X1 port map( A => n77, B => n90, S => A(21), Z => n67);
   U98 : MUX2_X1 port map( A => n88, B => n84, S => A(22), Z => n66);
   U99 : NAND3_X1 port map( A1 => n67, A2 => n86, A3 => n66, ZN => p_22_port);
   U100 : MUX2_X1 port map( A => n77, B => n90, S => A(22), Z => n69);
   U101 : MUX2_X1 port map( A => n88, B => n84, S => A(23), Z => n68);
   U102 : NAND3_X1 port map( A1 => n69, A2 => n86, A3 => n68, ZN => p_23_port);
   U103 : MUX2_X1 port map( A => n78, B => n90, S => A(23), Z => n71);
   U105 : NAND3_X1 port map( A1 => n71, A2 => n86, A3 => n88, ZN => p_24_port);
   U108 : NAND3_X1 port map( A1 => n77, A2 => n86, A3 => n88, ZN => p_25_port);
   U111 : NAND3_X1 port map( A1 => n78, A2 => n86, A3 => n88, ZN => p_26_port);
   U117 : NAND3_X1 port map( A1 => n78, A2 => n86, A3 => n88, ZN => p_28_port);
   U120 : NAND3_X1 port map( A1 => n78, A2 => n86, A3 => n88, ZN => p_29_port);
   U9 : NAND2_X1 port map( A1 => n17, A2 => b(2), ZN => n73);
   U10 : OR2_X2 port map( A1 => n19, A2 => b(2), ZN => n84);
   U8 : NAND2_X1 port map( A1 => b(1), A2 => b(0), ZN => n90);
   U5 : NAND2_X2 port map( A1 => b(2), A2 => n23, ZN => n86);
   U3 : OR2_X1 port map( A1 => n73, A2 => b(0), ZN => n78);
   U4 : OR2_X1 port map( A1 => n73, A2 => b(0), ZN => n77);
   U11 : INV_X1 port map( A => b(1), ZN => n17);
   U12 : OR2_X1 port map( A1 => n73, A2 => b(0), ZN => n89);
   U6 : OAI21_X2 port map( B1 => b(0), B2 => b(1), A => b(2), ZN => n88);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_9 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_9;

architecture SYN_beh of ENC_9 is

   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n6, n19, n20, n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, 
      n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47
      , n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
      n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n74, n87, n89, n91
      , n92, n93, n97, n98, n101 : std_logic;

begin
   
   U7 : AND2_X1 port map( A1 => n25, A2 => n26, ZN => n1);
   U12 : NAND3_X1 port map( A1 => n87, A2 => n93, A3 => n1, ZN => n89);
   U20 : XNOR2_X1 port map( A => b(0), B => b(1), ZN => n19);
   U25 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n21);
   U29 : NAND2_X1 port map( A1 => b(2), A2 => n21, ZN => n25);
   U30 : MUX2_X1 port map( A => n25, B => n87, S => A(0), Z => n20);
   U31 : OAI211_X1 port map( C1 => n22, C2 => n21, A => n92, B => n20, ZN => 
                           p(0));
   U33 : MUX2_X1 port map( A => n92, B => n93, S => A(0), Z => n28);
   U36 : MUX2_X1 port map( A => n91, B => n87, S => A(1), Z => n27);
   U37 : NAND3_X1 port map( A1 => n28, A2 => n101, A3 => n27, ZN => p(1));
   U38 : MUX2_X1 port map( A => n92, B => n93, S => A(1), Z => n30);
   U39 : MUX2_X1 port map( A => n91, B => n87, S => A(2), Z => n29);
   U40 : NAND3_X1 port map( A1 => n30, A2 => n6, A3 => n29, ZN => p(2));
   U41 : MUX2_X1 port map( A => n92, B => n93, S => A(2), Z => n32);
   U42 : MUX2_X1 port map( A => n91, B => n87, S => A(3), Z => n31);
   U43 : NAND3_X1 port map( A1 => n32, A2 => n101, A3 => n31, ZN => p(3));
   U44 : MUX2_X1 port map( A => n92, B => n93, S => A(3), Z => n34);
   U45 : MUX2_X1 port map( A => n91, B => n87, S => A(4), Z => n33);
   U46 : NAND3_X1 port map( A1 => n34, A2 => n6, A3 => n33, ZN => p(4));
   U47 : MUX2_X1 port map( A => n92, B => n93, S => A(4), Z => n36);
   U48 : MUX2_X1 port map( A => n91, B => n87, S => A(5), Z => n35);
   U49 : NAND3_X1 port map( A1 => n36, A2 => n101, A3 => n35, ZN => p(5));
   U50 : MUX2_X1 port map( A => n92, B => n93, S => A(5), Z => n38);
   U51 : MUX2_X1 port map( A => n91, B => n87, S => A(6), Z => n37);
   U52 : NAND3_X1 port map( A1 => n38, A2 => n6, A3 => n37, ZN => p(6));
   U53 : MUX2_X1 port map( A => n92, B => n93, S => A(6), Z => n40);
   U54 : MUX2_X1 port map( A => n91, B => n87, S => A(7), Z => n39);
   U55 : NAND3_X1 port map( A1 => n40, A2 => n6, A3 => n39, ZN => p(7));
   U56 : MUX2_X1 port map( A => n92, B => n93, S => A(7), Z => n42);
   U57 : MUX2_X1 port map( A => n91, B => n87, S => A(8), Z => n41);
   U58 : NAND3_X1 port map( A1 => n42, A2 => n101, A3 => n41, ZN => p(8));
   U59 : MUX2_X1 port map( A => n92, B => n93, S => A(8), Z => n44);
   U60 : MUX2_X1 port map( A => n91, B => n87, S => A(9), Z => n43);
   U61 : NAND3_X1 port map( A1 => n44, A2 => n6, A3 => n43, ZN => p(9));
   U62 : MUX2_X1 port map( A => n91, B => n87, S => A(10), Z => n46);
   U63 : MUX2_X1 port map( A => n92, B => n93, S => A(9), Z => n45);
   U64 : NAND3_X1 port map( A1 => n46, A2 => n101, A3 => n45, ZN => p(10));
   U65 : MUX2_X1 port map( A => n92, B => n93, S => A(10), Z => n48);
   U66 : MUX2_X1 port map( A => n91, B => n87, S => A(11), Z => n47);
   U67 : NAND3_X1 port map( A1 => n48, A2 => n101, A3 => n47, ZN => p(11));
   U68 : MUX2_X1 port map( A => n92, B => n93, S => A(11), Z => n50);
   U69 : MUX2_X1 port map( A => n91, B => n87, S => A(12), Z => n49);
   U70 : NAND3_X1 port map( A1 => n50, A2 => n101, A3 => n49, ZN => p(12));
   U71 : MUX2_X1 port map( A => n91, B => n87, S => A(13), Z => n52);
   U72 : MUX2_X1 port map( A => n92, B => n93, S => A(12), Z => n51);
   U73 : NAND3_X1 port map( A1 => n52, A2 => n101, A3 => n51, ZN => p(13));
   U74 : MUX2_X1 port map( A => n91, B => n87, S => A(14), Z => n54);
   U75 : MUX2_X1 port map( A => n92, B => n93, S => A(13), Z => n53);
   U76 : NAND3_X1 port map( A1 => n101, A2 => n54, A3 => n53, ZN => p(14));
   U77 : MUX2_X1 port map( A => n91, B => n87, S => A(15), Z => n56);
   U78 : MUX2_X1 port map( A => n92, B => n93, S => A(14), Z => n55);
   U79 : NAND3_X1 port map( A1 => n56, A2 => n6, A3 => n55, ZN => p(15));
   U80 : MUX2_X1 port map( A => n92, B => n93, S => A(15), Z => n58);
   U81 : MUX2_X1 port map( A => n91, B => n87, S => A(16), Z => n57);
   U82 : NAND3_X1 port map( A1 => n58, A2 => n6, A3 => n57, ZN => p(16));
   U83 : MUX2_X1 port map( A => n92, B => n93, S => A(16), Z => n60);
   U84 : MUX2_X1 port map( A => n91, B => n87, S => A(17), Z => n59);
   U85 : NAND3_X1 port map( A1 => n60, A2 => n6, A3 => n59, ZN => p(17));
   U86 : MUX2_X1 port map( A => n92, B => n93, S => A(17), Z => n62);
   U87 : MUX2_X1 port map( A => n91, B => n87, S => A(18), Z => n61);
   U88 : NAND3_X1 port map( A1 => n62, A2 => n101, A3 => n61, ZN => p(18));
   U89 : MUX2_X1 port map( A => n91, B => n87, S => A(19), Z => n64);
   U90 : MUX2_X1 port map( A => n92, B => n93, S => A(18), Z => n63);
   U91 : NAND3_X1 port map( A1 => n64, A2 => n63, A3 => n6, ZN => p(19));
   U92 : MUX2_X1 port map( A => n92, B => n93, S => A(19), Z => n66);
   U93 : MUX2_X1 port map( A => n91, B => n87, S => A(20), Z => n65);
   U94 : NAND3_X1 port map( A1 => n66, A2 => n101, A3 => n65, ZN => p(20));
   U95 : MUX2_X1 port map( A => n92, B => n93, S => A(20), Z => n68);
   U96 : MUX2_X1 port map( A => n91, B => n87, S => A(21), Z => n67);
   U97 : NAND3_X1 port map( A1 => n68, A2 => n101, A3 => n67, ZN => p(21));
   U98 : MUX2_X1 port map( A => n91, B => n87, S => A(22), Z => n70);
   U99 : MUX2_X1 port map( A => n92, B => n93, S => A(21), Z => n69);
   U100 : NAND3_X1 port map( A1 => n70, A2 => n101, A3 => n69, ZN => p(22));
   U101 : MUX2_X1 port map( A => n92, B => n93, S => A(22), Z => n72);
   U102 : MUX2_X1 port map( A => n91, B => n87, S => A(23), Z => n71);
   U103 : NAND3_X1 port map( A1 => n72, A2 => n101, A3 => n71, ZN => p(23));
   U104 : MUX2_X1 port map( A => n92, B => n93, S => A(23), Z => n74);
   U106 : NAND3_X1 port map( A1 => n74, A2 => n6, A3 => n91, ZN => p(24));
   U109 : NAND3_X1 port map( A1 => n92, A2 => n6, A3 => n91, ZN => p(25));
   U112 : NAND3_X1 port map( A1 => n92, A2 => n101, A3 => n91, ZN => p(26));
   U115 : NAND3_X1 port map( A1 => n92, A2 => n101, A3 => n91, ZN => p(27));
   U118 : NAND3_X1 port map( A1 => n92, A2 => n101, A3 => n91, ZN => p(28));
   U121 : NAND3_X1 port map( A1 => n92, A2 => n6, A3 => n91, ZN => p(29));
   U124 : NAND3_X1 port map( A1 => n92, A2 => n6, A3 => n91, ZN => p(30));
   U127 : NAND3_X1 port map( A1 => n92, A2 => n6, A3 => n91, ZN => p(31));
   U8 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n26);
   U9 : INV_X1 port map( A => b(0), ZN => n98);
   U16 : NAND3_X2 port map( A1 => n98, A2 => n97, A3 => b(2), ZN => n92);
   U3 : CLKBUF_X2 port map( A => n89, Z => n6);
   U35 : NAND2_X2 port map( A1 => b(2), A2 => n26, ZN => n91);
   U32 : NAND3_X1 port map( A1 => b(1), A2 => n22, A3 => b(0), ZN => n93);
   U4 : CLKBUF_X3 port map( A => n89, Z => n101);
   U5 : INV_X1 port map( A => b(1), ZN => n97);
   U10 : INV_X1 port map( A => b(2), ZN => n22);
   U6 : OR2_X2 port map( A1 => n19, A2 => b(2), ZN => n87);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_10 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_10;

architecture SYN_beh of ENC_10 is

   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal p_32_port, p_30_port, p_31_port, p_28_port, p_26_port, p_25_port, 
      p_24_port, p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, 
      p_18_port, p_17_port, p_16_port, p_15_port, p_14_port, p_13_port, 
      p_12_port, p_11_port, p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, 
      p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, p_0_port, n1, n3, n4, 
      n5, n6, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, n56, n57, n58, n59, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n75, n76, n78, n80, n89, n91, n93, n94
      , n96, n100, n101, n102, n103, n104 : std_logic;

begin
   p <= ( p_32_port, p_31_port, p_30_port, p_31_port, p_28_port, p_28_port, 
      p_26_port, p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, 
      p_20_port, p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, 
      p_14_port, p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port
      , p_7_port, p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, 
      p_0_port );
   
   U8 : NAND2_X1 port map( A1 => b(0), A2 => n100, ZN => n3);
   U9 : NAND2_X1 port map( A1 => n1, A2 => b(1), ZN => n4);
   U10 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n6);
   U11 : INV_X1 port map( A => b(0), ZN => n1);
   U24 : NAND3_X1 port map( A1 => b(1), A2 => b(0), A3 => b(2), ZN => n24);
   U27 : NAND2_X1 port map( A1 => n5, A2 => n100, ZN => n94);
   U30 : MUX2_X1 port map( A => n43, B => n89, S => A(0), Z => n23);
   U31 : NAND3_X1 port map( A1 => n24, A2 => n94, A3 => n23, ZN => p_0_port);
   U33 : MUX2_X1 port map( A => n94, B => n93, S => A(0), Z => n26);
   U36 : MUX2_X1 port map( A => n104, B => n89, S => A(1), Z => n25);
   U37 : NAND3_X1 port map( A1 => n26, A2 => n91, A3 => n25, ZN => p_1_port);
   U38 : MUX2_X1 port map( A => n78, B => n93, S => A(1), Z => n28);
   U39 : MUX2_X1 port map( A => n104, B => n102, S => A(2), Z => n27);
   U40 : NAND3_X1 port map( A1 => n28, A2 => n91, A3 => n27, ZN => p_2_port);
   U41 : MUX2_X1 port map( A => n94, B => n93, S => A(2), Z => n30);
   U42 : MUX2_X1 port map( A => n104, B => n101, S => A(3), Z => n29);
   U43 : NAND3_X1 port map( A1 => n30, A2 => n91, A3 => n29, ZN => p_3_port);
   U44 : MUX2_X1 port map( A => n94, B => n93, S => A(3), Z => n32);
   U45 : MUX2_X1 port map( A => n104, B => n89, S => A(4), Z => n31);
   U46 : NAND3_X1 port map( A1 => n32, A2 => n91, A3 => n31, ZN => p_4_port);
   U47 : MUX2_X1 port map( A => n94, B => n93, S => A(4), Z => n34);
   U48 : MUX2_X1 port map( A => n104, B => n102, S => A(5), Z => n33);
   U49 : NAND3_X1 port map( A1 => n34, A2 => n91, A3 => n33, ZN => p_5_port);
   U50 : MUX2_X1 port map( A => n94, B => n93, S => A(5), Z => n36);
   U51 : MUX2_X1 port map( A => n104, B => n89, S => A(6), Z => n35);
   U52 : NAND3_X1 port map( A1 => n36, A2 => n91, A3 => n35, ZN => p_6_port);
   U53 : MUX2_X1 port map( A => n78, B => n93, S => A(6), Z => n38);
   U54 : MUX2_X1 port map( A => n104, B => n101, S => A(7), Z => n37);
   U55 : NAND3_X1 port map( A1 => n38, A2 => n91, A3 => n37, ZN => p_7_port);
   U56 : MUX2_X1 port map( A => n104, B => n89, S => A(8), Z => n40);
   U57 : MUX2_X1 port map( A => n94, B => n93, S => A(7), Z => n39);
   U58 : NAND3_X1 port map( A1 => n40, A2 => n91, A3 => n39, ZN => p_8_port);
   U59 : MUX2_X1 port map( A => n78, B => n93, S => A(8), Z => n42);
   U60 : MUX2_X1 port map( A => n104, B => n89, S => A(9), Z => n41);
   U61 : NAND3_X1 port map( A1 => n42, A2 => n91, A3 => n41, ZN => p_9_port);
   U62 : MUX2_X1 port map( A => n94, B => n93, S => A(9), Z => n45);
   U63 : NAND2_X1 port map( A1 => n6, A2 => n43, ZN => n76);
   U64 : MUX2_X1 port map( A => n104, B => n89, S => A(10), Z => n44);
   U65 : NAND3_X1 port map( A1 => n45, A2 => n91, A3 => n44, ZN => p_10_port);
   U66 : MUX2_X1 port map( A => n78, B => n93, S => A(10), Z => n47);
   U67 : MUX2_X1 port map( A => n104, B => n89, S => A(11), Z => n46);
   U68 : NAND3_X1 port map( A1 => n47, A2 => n91, A3 => n46, ZN => p_11_port);
   U69 : MUX2_X1 port map( A => n78, B => n93, S => A(11), Z => n49);
   U70 : MUX2_X1 port map( A => n104, B => n102, S => A(12), Z => n48);
   U71 : NAND3_X1 port map( A1 => n49, A2 => n91, A3 => n48, ZN => p_12_port);
   U72 : MUX2_X1 port map( A => n78, B => n93, S => A(12), Z => n51);
   U73 : MUX2_X1 port map( A => n104, B => n89, S => A(13), Z => n50);
   U74 : NAND3_X1 port map( A1 => n51, A2 => n91, A3 => n50, ZN => p_13_port);
   U75 : MUX2_X1 port map( A => n78, B => n93, S => A(13), Z => n53);
   U76 : MUX2_X1 port map( A => n96, B => n76, S => A(14), Z => n52);
   U77 : NAND3_X1 port map( A1 => n53, A2 => n91, A3 => n52, ZN => p_14_port);
   U78 : MUX2_X1 port map( A => n78, B => n93, S => A(14), Z => n55);
   U79 : MUX2_X1 port map( A => n96, B => n76, S => A(15), Z => n54);
   U80 : NAND3_X1 port map( A1 => n55, A2 => n91, A3 => n54, ZN => p_15_port);
   U81 : MUX2_X1 port map( A => n78, B => n93, S => A(15), Z => n57);
   U82 : MUX2_X1 port map( A => n96, B => n76, S => A(16), Z => n56);
   U83 : NAND3_X1 port map( A1 => n57, A2 => n91, A3 => n56, ZN => p_16_port);
   U84 : MUX2_X1 port map( A => n96, B => n76, S => A(17), Z => n59);
   U85 : MUX2_X1 port map( A => n94, B => n93, S => A(16), Z => n58);
   U86 : NAND3_X1 port map( A1 => n91, A2 => n59, A3 => n58, ZN => p_17_port);
   U87 : NAND2_X1 port map( A1 => n5, A2 => n100, ZN => n78);
   U88 : MUX2_X1 port map( A => n94, B => n93, S => A(17), Z => n63);
   U89 : MUX2_X1 port map( A => n96, B => n101, S => A(18), Z => n62);
   U90 : NAND3_X1 port map( A1 => n63, A2 => n91, A3 => n62, ZN => p_18_port);
   U91 : MUX2_X1 port map( A => n78, B => n93, S => A(18), Z => n65);
   U92 : MUX2_X1 port map( A => n104, B => n102, S => A(19), Z => n64);
   U93 : NAND3_X1 port map( A1 => n65, A2 => n91, A3 => n64, ZN => p_19_port);
   U94 : MUX2_X1 port map( A => n94, B => n93, S => A(19), Z => n67);
   U95 : MUX2_X1 port map( A => n104, B => n89, S => A(20), Z => n66);
   U96 : NAND3_X1 port map( A1 => n67, A2 => n91, A3 => n66, ZN => p_20_port);
   U97 : MUX2_X1 port map( A => n104, B => n89, S => A(21), Z => n69);
   U98 : MUX2_X1 port map( A => n80, B => n93, S => A(20), Z => n68);
   U99 : NAND3_X1 port map( A1 => n69, A2 => n91, A3 => n68, ZN => p_21_port);
   U100 : MUX2_X1 port map( A => n80, B => n93, S => A(21), Z => n71);
   U101 : MUX2_X1 port map( A => n104, B => n102, S => A(22), Z => n70);
   U102 : NAND3_X1 port map( A1 => n71, A2 => n91, A3 => n70, ZN => p_22_port);
   U103 : MUX2_X1 port map( A => n80, B => n93, S => A(22), Z => n73);
   U104 : MUX2_X1 port map( A => n104, B => n102, S => A(23), Z => n72);
   U105 : NAND3_X1 port map( A1 => n72, A2 => n91, A3 => n73, ZN => p_23_port);
   U106 : MUX2_X1 port map( A => n80, B => n93, S => A(23), Z => n75);
   U108 : NAND3_X1 port map( A1 => n75, A2 => n91, A3 => n104, ZN => p_24_port)
                           ;
   U111 : NAND3_X1 port map( A1 => n78, A2 => n91, A3 => n104, ZN => p_25_port)
                           ;
   U114 : NAND3_X1 port map( A1 => n80, A2 => n91, A3 => n104, ZN => p_26_port)
                           ;
   U117 : NAND3_X1 port map( A1 => n80, A2 => n91, A3 => n104, ZN => p_28_port)
                           ;
   U123 : NAND3_X1 port map( A1 => n80, A2 => n91, A3 => n104, ZN => p_31_port)
                           ;
   U126 : NAND3_X1 port map( A1 => n80, A2 => n91, A3 => n104, ZN => p_30_port)
                           ;
   U131 : NAND2_X1 port map( A1 => n104, A2 => n80, ZN => p_32_port);
   U3 : NAND2_X1 port map( A1 => n100, A2 => n5, ZN => n80);
   U5 : AND2_X1 port map( A1 => b(2), A2 => n1, ZN => n5);
   U7 : NAND2_X1 port map( A1 => n103, A2 => n43, ZN => n101);
   U13 : NAND2_X1 port map( A1 => n103, A2 => n43, ZN => n102);
   U16 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => n103);
   U17 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n93);
   U19 : NAND2_X1 port map( A1 => n103, A2 => n43, ZN => n89);
   U20 : INV_X1 port map( A => b(1), ZN => n100);
   U15 : BUF_X1 port map( A => n96, Z => n104);
   U4 : INV_X1 port map( A => b(2), ZN => n43);
   U6 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => b(2), ZN => n96);
   U12 : NAND3_X2 port map( A1 => b(0), A2 => b(2), A3 => b(1), ZN => n91);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_11 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_11;

architecture SYN_beh of ENC_11 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal p_32_port, p_31_port, p_30_port, p_29_port, p_27_port, p_26_port, 
      p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, p_20_port, 
      p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, p_14_port, 
      p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port, p_7_port,
      p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, p_0_port, n1,
      n2, n5, n7, n9, n10, n15, n17, n18, n19, n27, n28, n32, n34, n35, n36, 
      n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52
      , n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n93, n97, n98, n99, 
      n102, n107, n116, n119, n120, n121, n122 : std_logic;

begin
   p <= ( p_32_port, p_31_port, p_30_port, p_29_port, p_30_port, p_27_port, 
      p_26_port, p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, 
      p_20_port, p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, 
      p_14_port, p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port
      , p_7_port, p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, 
      p_0_port );
   
   U3 : NAND2_X1 port map( A1 => A(21), A2 => n15, ZN => n1);
   U4 : NAND2_X1 port map( A1 => n32, A2 => n34, ZN => n2);
   U5 : AND3_X1 port map( A1 => n1, A2 => n2, A3 => n17, ZN => n86);
   U6 : NAND3_X1 port map( A1 => n17, A2 => n58, A3 => n59, ZN => p_11_port);
   U12 : NAND2_X1 port map( A1 => n7, A2 => n79, ZN => n5);
   U15 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n7);
   U17 : NAND2_X1 port map( A1 => b(0), A2 => n116, ZN => n9);
   U19 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n19);
   U26 : INV_X1 port map( A => n97, ZN => n15);
   U37 : INV_X1 port map( A => n98, ZN => n32);
   U39 : INV_X1 port map( A => A(21), ZN => n34);
   U42 : INV_X1 port map( A => b(0), ZN => n35);
   U44 : NAND2_X1 port map( A1 => b(2), A2 => n73, ZN => n72);
   U45 : NAND2_X1 port map( A1 => n19, A2 => n79, ZN => n107);
   U46 : MUX2_X1 port map( A => n72, B => n97, S => A(0), Z => n36);
   U47 : OAI211_X1 port map( C1 => n79, C2 => n28, A => n99, B => n36, ZN => 
                           p_0_port);
   U48 : MUX2_X1 port map( A => n99, B => n28, S => A(0), Z => n39);
   U51 : OAI21_X1 port map( B1 => b(0), B2 => b(1), A => b(2), ZN => n98);
   U53 : NAND3_X1 port map( A1 => n39, A2 => n17, A3 => n38, ZN => p_1_port);
   U54 : MUX2_X1 port map( A => n122, B => n28, S => A(1), Z => n41);
   U56 : NAND3_X1 port map( A1 => n41, A2 => n17, A3 => n40, ZN => p_2_port);
   U57 : MUX2_X1 port map( A => n102, B => n28, S => A(2), Z => n43);
   U59 : NAND3_X1 port map( A1 => n43, A2 => n17, A3 => n42, ZN => p_3_port);
   U60 : MUX2_X1 port map( A => n102, B => n28, S => A(3), Z => n45);
   U62 : NAND3_X1 port map( A1 => n45, A2 => n17, A3 => n44, ZN => p_4_port);
   U65 : NAND3_X1 port map( A1 => n47, A2 => n17, A3 => n46, ZN => p_5_port);
   U66 : MUX2_X1 port map( A => n99, B => n28, S => A(5), Z => n49);
   U68 : NAND3_X1 port map( A1 => n49, A2 => n17, A3 => n48, ZN => p_6_port);
   U71 : NAND3_X1 port map( A1 => n51, A2 => n17, A3 => n50, ZN => p_7_port);
   U72 : MUX2_X1 port map( A => n99, B => n28, S => A(7), Z => n53);
   U74 : NAND3_X1 port map( A1 => n53, A2 => n17, A3 => n52, ZN => p_8_port);
   U75 : MUX2_X1 port map( A => n122, B => n28, S => A(8), Z => n55);
   U77 : NAND3_X1 port map( A1 => n55, A2 => n17, A3 => n54, ZN => p_9_port);
   U79 : MUX2_X1 port map( A => n102, B => n27, S => A(9), Z => n56);
   U80 : NAND3_X1 port map( A1 => n57, A2 => n17, A3 => n56, ZN => p_10_port);
   U81 : MUX2_X1 port map( A => n99, B => n27, S => A(10), Z => n59);
   U83 : MUX2_X1 port map( A => n122, B => n27, S => A(11), Z => n61);
   U85 : NAND3_X1 port map( A1 => n61, A2 => n17, A3 => n60, ZN => p_12_port);
   U86 : MUX2_X1 port map( A => n102, B => n27, S => A(12), Z => n63);
   U88 : NAND3_X1 port map( A1 => n63, A2 => n17, A3 => n62, ZN => p_13_port);
   U89 : MUX2_X1 port map( A => n99, B => n27, S => A(13), Z => n65);
   U91 : NAND3_X1 port map( A1 => n65, A2 => n17, A3 => n64, ZN => p_14_port);
   U92 : MUX2_X1 port map( A => n99, B => n27, S => A(14), Z => n67);
   U94 : NAND3_X1 port map( A1 => n67, A2 => n17, A3 => n66, ZN => p_15_port);
   U95 : MUX2_X1 port map( A => n99, B => n27, S => A(15), Z => n69);
   U96 : NAND2_X1 port map( A1 => n19, A2 => n79, ZN => n97);
   U97 : MUX2_X1 port map( A => n82, B => n5, S => A(16), Z => n68);
   U98 : NAND3_X1 port map( A1 => n69, A2 => n17, A3 => n68, ZN => p_16_port);
   U99 : MUX2_X1 port map( A => n122, B => n27, S => A(16), Z => n71);
   U100 : MUX2_X1 port map( A => n93, B => n5, S => A(17), Z => n70);
   U101 : NAND3_X1 port map( A1 => n71, A2 => n17, A3 => n70, ZN => p_17_port);
   U102 : INV_X1 port map( A => n72, ZN => n76);
   U104 : MUX2_X1 port map( A => n82, B => n107, S => A(18), Z => n74);
   U105 : OAI211_X1 port map( C1 => n76, C2 => n93, A => n74, B => n75, ZN => 
                           p_18_port);
   U106 : MUX2_X1 port map( A => n82, B => n97, S => A(19), Z => n78);
   U107 : MUX2_X1 port map( A => n120, B => n27, S => A(18), Z => n77);
   U108 : NAND3_X1 port map( A1 => n17, A2 => n78, A3 => n77, ZN => p_19_port);
   U109 : XOR2_X1 port map( A => b(1), B => b(0), Z => n80);
   U110 : NAND2_X1 port map( A1 => n80, A2 => n79, ZN => n81);
   U111 : MUX2_X1 port map( A => n82, B => n81, S => A(20), Z => n84);
   U112 : MUX2_X1 port map( A => n99, B => n27, S => A(19), Z => n83);
   U113 : NAND3_X1 port map( A1 => n84, A2 => n17, A3 => n83, ZN => p_20_port);
   U114 : MUX2_X1 port map( A => n99, B => n27, S => A(20), Z => n85);
   U115 : NAND2_X1 port map( A1 => n86, A2 => n85, ZN => p_21_port);
   U116 : MUX2_X1 port map( A => n102, B => n28, S => A(21), Z => n88);
   U117 : MUX2_X1 port map( A => n93, B => n5, S => A(22), Z => n87);
   U118 : NAND3_X1 port map( A1 => n88, A2 => n17, A3 => n87, ZN => p_22_port);
   U120 : MUX2_X1 port map( A => n122, B => n28, S => A(22), Z => n89);
   U121 : NAND3_X1 port map( A1 => n90, A2 => n17, A3 => n89, ZN => p_23_port);
   U124 : NAND3_X1 port map( A1 => n92, A2 => n17, A3 => n93, ZN => p_24_port);
   U130 : NAND3_X1 port map( A1 => n98, A2 => n17, A3 => n102, ZN => p_26_port)
                           ;
   U136 : NAND3_X1 port map( A1 => n122, A2 => n17, A3 => n98, ZN => p_27_port)
                           ;
   U139 : NAND3_X1 port map( A1 => n122, A2 => n93, A3 => n17, ZN => p_29_port)
                           ;
   U142 : NAND3_X1 port map( A1 => n99, A2 => n17, A3 => n98, ZN => p_30_port);
   U147 : NAND2_X1 port map( A1 => n98, A2 => n102, ZN => p_32_port);
   U10 : NAND2_X1 port map( A1 => n18, A2 => n116, ZN => n102);
   U11 : NAND2_X1 port map( A1 => n18, A2 => n116, ZN => n120);
   U13 : AND2_X1 port map( A1 => n93, A2 => n120, ZN => n119);
   U18 : NAND2_X1 port map( A1 => n17, A2 => n119, ZN => p_25_port);
   U20 : OAI21_X1 port map( B1 => b(1), B2 => b(0), A => b(2), ZN => n82);
   U21 : MUX2_X1 port map( A => n120, B => n73, S => A(17), Z => n75);
   U22 : MUX2_X1 port map( A => n122, B => n28, S => A(23), Z => n92);
   U23 : MUX2_X1 port map( A => n122, B => n28, S => A(4), Z => n47);
   U25 : MUX2_X1 port map( A => n102, B => n28, S => A(6), Z => n51);
   U29 : NAND2_X1 port map( A1 => n17, A2 => n119, ZN => p_31_port);
   U30 : MUX2_X1 port map( A => n98, B => n121, S => A(3), Z => n42);
   U31 : MUX2_X1 port map( A => n98, B => n121, S => A(23), Z => n90);
   U32 : MUX2_X1 port map( A => n93, B => n121, S => A(12), Z => n60);
   U34 : MUX2_X1 port map( A => n93, B => n121, S => A(11), Z => n58);
   U35 : MUX2_X1 port map( A => n98, B => n121, S => A(14), Z => n64);
   U38 : MUX2_X1 port map( A => n93, B => n121, S => A(8), Z => n52);
   U49 : MUX2_X1 port map( A => n93, B => n121, S => A(5), Z => n46);
   U50 : MUX2_X1 port map( A => n93, B => n121, S => A(10), Z => n57);
   U52 : MUX2_X1 port map( A => n93, B => n121, S => A(6), Z => n48);
   U55 : MUX2_X1 port map( A => n98, B => n121, S => A(9), Z => n54);
   U58 : MUX2_X1 port map( A => n93, B => n121, S => A(15), Z => n66);
   U61 : MUX2_X1 port map( A => n98, B => n121, S => A(4), Z => n44);
   U63 : MUX2_X1 port map( A => n98, B => n121, S => A(2), Z => n40);
   U64 : MUX2_X1 port map( A => n98, B => n121, S => A(7), Z => n50);
   U67 : MUX2_X1 port map( A => n93, B => n121, S => A(1), Z => n38);
   U69 : MUX2_X1 port map( A => n93, B => n121, S => A(13), Z => n62);
   U76 : OR2_X1 port map( A1 => b(0), A2 => n116, ZN => n10);
   U78 : NAND2_X1 port map( A1 => n18, A2 => n116, ZN => n122);
   U33 : AND2_X1 port map( A1 => b(2), A2 => n35, ZN => n18);
   U14 : CLKBUF_X1 port map( A => n73, Z => n27);
   U43 : NAND2_X1 port map( A1 => n18, A2 => n116, ZN => n99);
   U70 : NAND2_X1 port map( A1 => n7, A2 => n79, ZN => n121);
   U41 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n73);
   U16 : CLKBUF_X1 port map( A => n73, Z => n28);
   U8 : NAND2_X4 port map( A1 => n32, A2 => n72, ZN => n17);
   U9 : INV_X1 port map( A => b(1), ZN => n116);
   U27 : INV_X1 port map( A => b(2), ZN => n79);
   U7 : INV_X2 port map( A => n32, ZN => n93);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_12 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_12;

architecture SYN_beh of ENC_12 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net29919, net29922, net29924, net29930, net29949, net31213, net31510,
      net31509, net31508, net29996, net29995, net29994, net29951, net29948, 
      net29921, net37587, net34501, net29964, net34125, net29926, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n79, n80, n81, n82, n83 : std_logic;

begin
   
   U7 : NAND2_X1 port map( A1 => net29964, A2 => n5, ZN => net31213);
   U8 : NAND2_X1 port map( A1 => net34125, A2 => b(2), ZN => net29926);
   U10 : NAND2_X1 port map( A1 => b(2), A2 => net34125, ZN => net29919);
   U14 : NAND2_X1 port map( A1 => net31508, A2 => n67, ZN => net34125);
   U17 : NAND2_X1 port map( A1 => b(2), A2 => net29995, ZN => net29994);
   U18 : INV_X1 port map( A => b(2), ZN => net29964);
   U20 : NAND2_X1 port map( A1 => net37587, A2 => net29964, ZN => net34501);
   U22 : NAND2_X1 port map( A1 => n5, A2 => net29964, ZN => net29930);
   U23 : OAI211_X1 port map( C1 => net29964, C2 => net29922, A => net29921, B 
                           => net29996, ZN => p(0));
   U25 : NAND2_X1 port map( A1 => net31509, A2 => net31510, ZN => n5);
   U26 : MUX2_X1 port map( A => net29921, B => net29922, S => A(19), Z => 
                           net29949);
   U29 : NAND3_X1 port map( A1 => net29948, A2 => n6, A3 => net29924, ZN => 
                           p(21));
   U30 : MUX2_X1 port map( A => net29921, B => net29995, S => A(18), Z => 
                           net29951);
   U32 : MUX2_X1 port map( A => net29921, B => net29922, S => A(20), Z => n6);
   U33 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => net29995);
   U47 : NAND2_X1 port map( A1 => b(1), A2 => net31508, ZN => net31509);
   U48 : NAND2_X1 port map( A1 => b(0), A2 => n67, ZN => net31510);
   U50 : INV_X1 port map( A => b(0), ZN => net31508);
   U52 : MUX2_X1 port map( A => net29921, B => net29922, S => A(0), Z => n8);
   U54 : NAND3_X1 port map( A1 => n8, A2 => net29924, A3 => n7, ZN => p(1));
   U55 : MUX2_X1 port map( A => net29921, B => net29922, S => A(1), Z => n10);
   U57 : NAND3_X1 port map( A1 => n10, A2 => net29924, A3 => n9, ZN => p(2));
   U58 : MUX2_X1 port map( A => net29921, B => net29922, S => A(2), Z => n12);
   U60 : NAND3_X1 port map( A1 => n12, A2 => net29924, A3 => n11, ZN => p(3));
   U61 : MUX2_X1 port map( A => net29921, B => net29922, S => A(3), Z => n14);
   U63 : NAND3_X1 port map( A1 => n14, A2 => net29924, A3 => n13, ZN => p(4));
   U64 : MUX2_X1 port map( A => net29921, B => net29922, S => A(4), Z => n16);
   U66 : NAND3_X1 port map( A1 => n16, A2 => net29924, A3 => n15, ZN => p(5));
   U67 : MUX2_X1 port map( A => net29921, B => net29922, S => A(5), Z => n18);
   U68 : MUX2_X1 port map( A => n72, B => net31213, S => A(6), Z => n17);
   U69 : NAND3_X1 port map( A1 => n18, A2 => net29924, A3 => n17, ZN => p(6));
   U70 : MUX2_X1 port map( A => net29921, B => net29922, S => A(6), Z => n20);
   U71 : MUX2_X1 port map( A => n72, B => net31213, S => A(7), Z => n19);
   U72 : NAND3_X1 port map( A1 => n20, A2 => net29924, A3 => n19, ZN => p(7));
   U73 : MUX2_X1 port map( A => net29921, B => net29922, S => A(7), Z => n22);
   U74 : MUX2_X1 port map( A => n72, B => n83, S => A(8), Z => n21);
   U75 : NAND3_X1 port map( A1 => n22, A2 => net29924, A3 => n21, ZN => p(8));
   U76 : MUX2_X1 port map( A => net29921, B => net29922, S => A(8), Z => n24);
   U77 : MUX2_X1 port map( A => n72, B => net31213, S => A(9), Z => n23);
   U78 : NAND3_X1 port map( A1 => n24, A2 => net29924, A3 => n23, ZN => p(9));
   U79 : MUX2_X1 port map( A => net29921, B => net29922, S => A(9), Z => n26);
   U81 : NAND3_X1 port map( A1 => n26, A2 => net29924, A3 => n25, ZN => p(10));
   U82 : MUX2_X1 port map( A => net29921, B => net29922, S => A(10), Z => n28);
   U83 : MUX2_X1 port map( A => n72, B => n83, S => A(11), Z => n27);
   U84 : NAND3_X1 port map( A1 => n28, A2 => net29924, A3 => n27, ZN => p(11));
   U85 : MUX2_X1 port map( A => net29921, B => net29922, S => A(11), Z => n30);
   U87 : NAND3_X1 port map( A1 => n30, A2 => net29924, A3 => n29, ZN => p(12));
   U88 : MUX2_X1 port map( A => net29921, B => net29922, S => A(12), Z => n32);
   U89 : MUX2_X1 port map( A => n72, B => net29930, S => A(13), Z => n31);
   U90 : NAND3_X1 port map( A1 => n32, A2 => net29924, A3 => n31, ZN => p(13));
   U91 : MUX2_X1 port map( A => n47, B => net31213, S => A(14), Z => n34);
   U92 : MUX2_X1 port map( A => net29921, B => net29922, S => A(13), Z => n33);
   U93 : NAND3_X1 port map( A1 => n34, A2 => net29924, A3 => n33, ZN => p(14));
   U94 : MUX2_X1 port map( A => net29921, B => net29922, S => A(14), Z => n36);
   U95 : MUX2_X1 port map( A => n72, B => net31213, S => A(15), Z => n35);
   U96 : NAND3_X1 port map( A1 => n36, A2 => net29924, A3 => n35, ZN => p(15));
   U97 : MUX2_X1 port map( A => net29921, B => net29922, S => A(15), Z => n38);
   U99 : NAND3_X1 port map( A1 => n38, A2 => net29924, A3 => n37, ZN => p(16));
   U100 : MUX2_X1 port map( A => net29921, B => net29922, S => A(16), Z => n40)
                           ;
   U101 : MUX2_X1 port map( A => net29919, B => n83, S => A(17), Z => n39);
   U102 : NAND3_X1 port map( A1 => n40, A2 => net29924, A3 => n39, ZN => p(17))
                           ;
   U103 : MUX2_X1 port map( A => net29921, B => net29922, S => A(17), Z => n41)
                           ;
   U105 : MUX2_X1 port map( A => n72, B => net29930, S => A(20), Z => n42);
   U106 : NAND3_X1 port map( A1 => net29949, A2 => n42, A3 => net29924, ZN => 
                           p(20));
   U107 : MUX2_X1 port map( A => net29921, B => net29922, S => A(21), Z => n44)
                           ;
   U109 : NAND3_X1 port map( A1 => n44, A2 => net29924, A3 => n43, ZN => p(22))
                           ;
   U110 : MUX2_X1 port map( A => net29921, B => net29922, S => A(22), Z => n46)
                           ;
   U111 : MUX2_X1 port map( A => n72, B => n83, S => A(23), Z => n45);
   U112 : NAND3_X1 port map( A1 => n46, A2 => net29924, A3 => n45, ZN => p(23))
                           ;
   U113 : MUX2_X1 port map( A => net29921, B => net29922, S => A(23), Z => n48)
                           ;
   U115 : NAND3_X1 port map( A1 => n48, A2 => net29924, A3 => n47, ZN => p(24))
                           ;
   U118 : NAND3_X1 port map( A1 => net29921, A2 => net29924, A3 => net29919, ZN
                           => p(25));
   U121 : NAND3_X1 port map( A1 => net29921, A2 => net29924, A3 => net29919, ZN
                           => p(26));
   U124 : NAND3_X1 port map( A1 => net29921, A2 => net29924, A3 => n72, ZN => 
                           p(27));
   U127 : NAND3_X1 port map( A1 => net29921, A2 => net29924, A3 => n47, ZN => 
                           p(28));
   U130 : NAND3_X1 port map( A1 => net29921, A2 => net29924, A3 => n47, ZN => 
                           p(29));
   U133 : NAND3_X1 port map( A1 => net29921, A2 => net29924, A3 => net29919, ZN
                           => p(30));
   U136 : NAND3_X1 port map( A1 => net29921, A2 => net29924, A3 => n47, ZN => 
                           p(31));
   U138 : NAND2_X1 port map( A1 => n72, A2 => net29921, ZN => p(32));
   U3 : NAND3_X1 port map( A1 => net29951, A2 => n70, A3 => n68, ZN => p(19));
   U4 : INV_X1 port map( A => n69, ZN => n68);
   U9 : OAI21_X1 port map( B1 => net29926, B2 => A(19), A => net29924, ZN => 
                           n69);
   U16 : NAND2_X1 port map( A1 => b(2), A2 => net34125, ZN => n72);
   U24 : AOI21_X1 port map( B1 => n74, B2 => net29964, A => n75, ZN => n73);
   U27 : AND2_X1 port map( A1 => net37587, A2 => A(18), ZN => n74);
   U28 : AND3_X1 port map( A1 => net34125, A2 => b(2), A3 => n82, ZN => n75);
   U35 : NAND2_X1 port map( A1 => n5, A2 => net29964, ZN => n83);
   U39 : NAND2_X1 port map( A1 => net34125, A2 => b(2), ZN => n47);
   U43 : NAND2_X1 port map( A1 => net31509, A2 => net31510, ZN => net37587);
   U44 : INV_X1 port map( A => A(18), ZN => n82);
   U45 : NAND2_X1 port map( A1 => net34501, A2 => A(21), ZN => n81);
   U46 : NAND2_X1 port map( A1 => n81, A2 => n79, ZN => net29948);
   U49 : NAND2_X1 port map( A1 => net29919, A2 => n80, ZN => n79);
   U51 : INV_X1 port map( A => A(21), ZN => n80);
   U53 : NAND3_X1 port map( A1 => net29924, A2 => n41, A3 => n73, ZN => p(18));
   U56 : MUX2_X1 port map( A => n47, B => net29930, S => A(12), Z => n29);
   U59 : MUX2_X1 port map( A => n47, B => net29930, S => A(16), Z => n37);
   U62 : MUX2_X1 port map( A => n47, B => n83, S => A(22), Z => n43);
   U65 : MUX2_X1 port map( A => n47, B => n83, S => A(10), Z => n25);
   U80 : MUX2_X1 port map( A => net29994, B => n83, S => A(0), Z => net29996);
   U86 : MUX2_X1 port map( A => n72, B => n83, S => A(5), Z => n15);
   U98 : MUX2_X1 port map( A => n72, B => n83, S => A(4), Z => n13);
   U104 : MUX2_X1 port map( A => n72, B => n83, S => A(2), Z => n9);
   U108 : MUX2_X1 port map( A => net29919, B => n83, S => A(3), Z => n11);
   U114 : MUX2_X1 port map( A => n72, B => n83, S => A(1), Z => n7);
   U36 : NAND2_X2 port map( A1 => b(0), A2 => b(1), ZN => net29922);
   U13 : INV_X1 port map( A => A(19), ZN => n71);
   U15 : OR2_X1 port map( A1 => net34501, A2 => n71, ZN => n70);
   U19 : INV_X1 port map( A => b(1), ZN => n67);
   U5 : NAND3_X2 port map( A1 => net31508, A2 => b(2), A3 => n67, ZN => 
                           net29921);
   U6 : NAND2_X2 port map( A1 => net29994, A2 => b(2), ZN => net29924);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_13 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_13;

architecture SYN_beh of ENC_13 is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal p_32_port, p_31_port, p_30_port, p_29_port, p_27_port, p_26_port, 
      p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, p_20_port, 
      p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, p_14_port, 
      p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port, p_7_port,
      p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, p_0_port, 
      net29998, net30001, net30010, net30022, net30033, net30075, net30077, 
      net30721, net31233, net33597, net34028, net37654, net42472, net30030, 
      net33339, n1, n2, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n57, n58, n70, n72, n78
      , n83, n86, n87, n88 : std_logic;

begin
   p <= ( p_32_port, p_31_port, p_30_port, p_29_port, p_31_port, p_27_port, 
      p_26_port, p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, 
      p_20_port, p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, 
      p_14_port, p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port
      , p_7_port, p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, 
      p_0_port );
   
   U8 : INV_X1 port map( A => b(0), ZN => n1);
   U13 : NAND3_X1 port map( A1 => net30030, A2 => n2, A3 => net42472, ZN => 
                           p_21_port);
   U15 : MUX2_X1 port map( A => net30010, B => net29998, S => net30721, Z => n2
                           );
   U16 : NAND2_X1 port map( A1 => net33597, A2 => net30033, ZN => net30010);
   U18 : INV_X1 port map( A => A(21), ZN => net30721);
   U29 : INV_X1 port map( A => net29998, ZN => net37654);
   U31 : AND2_X1 port map( A1 => net37654, A2 => net30077, ZN => n5);
   U34 : AND2_X1 port map( A1 => net33339, A2 => net30721, ZN => n6);
   U35 : AND2_X1 port map( A1 => A(21), A2 => net31233, ZN => n7);
   U36 : NOR3_X1 port map( A1 => n5, A2 => n7, A3 => n6, ZN => n54);
   U37 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => net30075);
   U38 : XNOR2_X1 port map( A => b(0), B => n78, ZN => n8);
   U39 : XNOR2_X1 port map( A => b(0), B => n78, ZN => net33597);
   U40 : INV_X1 port map( A => net30001, ZN => net31233);
   U41 : NAND2_X1 port map( A1 => net33597, A2 => net30033, ZN => n9);
   U42 : INV_X1 port map( A => n5, ZN => n10);
   U44 : INV_X1 port map( A => b(2), ZN => net30033);
   U45 : NAND2_X1 port map( A1 => b(2), A2 => net30001, ZN => net30077);
   U46 : NAND2_X1 port map( A1 => n8, A2 => net30033, ZN => n70);
   U47 : MUX2_X1 port map( A => net30077, B => n70, S => A(0), Z => n11);
   U48 : OAI211_X1 port map( C1 => net30033, C2 => net30001, A => n88, B => n11
                           , ZN => p_0_port);
   U50 : MUX2_X1 port map( A => n88, B => net30001, S => A(0), Z => n13);
   U52 : MUX2_X1 port map( A => net29998, B => n70, S => A(1), Z => n12);
   U53 : NAND3_X1 port map( A1 => n13, A2 => n72, A3 => n12, ZN => p_1_port);
   U54 : MUX2_X1 port map( A => n88, B => net30001, S => A(1), Z => n15);
   U55 : MUX2_X1 port map( A => net29998, B => n70, S => A(2), Z => n14);
   U56 : NAND3_X1 port map( A1 => n15, A2 => n10, A3 => n14, ZN => p_2_port);
   U58 : MUX2_X1 port map( A => net29998, B => n70, S => A(3), Z => n16);
   U59 : NAND3_X1 port map( A1 => n17, A2 => n10, A3 => n16, ZN => p_3_port);
   U60 : MUX2_X1 port map( A => n88, B => net30001, S => A(3), Z => n19);
   U61 : MUX2_X1 port map( A => net29998, B => n70, S => A(4), Z => n18);
   U62 : NAND3_X1 port map( A1 => n19, A2 => n10, A3 => n18, ZN => p_4_port);
   U63 : MUX2_X1 port map( A => n88, B => net30001, S => A(4), Z => n21);
   U64 : MUX2_X1 port map( A => net29998, B => n9, S => A(5), Z => n20);
   U65 : NAND3_X1 port map( A1 => n21, A2 => n10, A3 => n20, ZN => p_5_port);
   U66 : MUX2_X1 port map( A => n88, B => net30001, S => A(5), Z => n23);
   U67 : MUX2_X1 port map( A => net29998, B => n70, S => A(6), Z => n22);
   U68 : NAND3_X1 port map( A1 => n23, A2 => n10, A3 => n22, ZN => p_6_port);
   U69 : MUX2_X1 port map( A => n88, B => net30001, S => A(6), Z => n25);
   U70 : MUX2_X1 port map( A => net29998, B => n9, S => A(7), Z => n24);
   U71 : NAND3_X1 port map( A1 => n25, A2 => n10, A3 => n24, ZN => p_7_port);
   U72 : MUX2_X1 port map( A => n88, B => net30001, S => A(7), Z => n27);
   U73 : MUX2_X1 port map( A => net29998, B => n70, S => A(8), Z => n26);
   U74 : NAND3_X1 port map( A1 => n27, A2 => n72, A3 => n26, ZN => p_8_port);
   U75 : MUX2_X1 port map( A => n88, B => net30001, S => A(8), Z => n29);
   U76 : MUX2_X1 port map( A => net29998, B => n70, S => A(9), Z => n28);
   U77 : NAND3_X1 port map( A1 => n29, A2 => net42472, A3 => n28, ZN => 
                           p_9_port);
   U78 : MUX2_X1 port map( A => n88, B => net30001, S => A(9), Z => n31);
   U79 : MUX2_X1 port map( A => n58, B => n9, S => A(10), Z => n30);
   U80 : NAND3_X1 port map( A1 => n31, A2 => net42472, A3 => n30, ZN => 
                           p_10_port);
   U81 : MUX2_X1 port map( A => n88, B => net30001, S => A(10), Z => n33);
   U82 : MUX2_X1 port map( A => n58, B => n70, S => A(11), Z => n32);
   U83 : NAND3_X1 port map( A1 => n33, A2 => net42472, A3 => n32, ZN => 
                           p_11_port);
   U84 : MUX2_X1 port map( A => n88, B => net30001, S => A(11), Z => n35);
   U85 : MUX2_X1 port map( A => n58, B => n9, S => A(12), Z => n34);
   U86 : NAND3_X1 port map( A1 => n35, A2 => net42472, A3 => n34, ZN => 
                           p_12_port);
   U87 : MUX2_X1 port map( A => n88, B => net30001, S => A(12), Z => n37);
   U88 : MUX2_X1 port map( A => n58, B => n70, S => A(13), Z => n36);
   U89 : NAND3_X1 port map( A1 => n37, A2 => n72, A3 => n36, ZN => p_13_port);
   U90 : MUX2_X1 port map( A => net29998, B => n9, S => A(14), Z => n39);
   U92 : NAND3_X1 port map( A1 => n39, A2 => n72, A3 => n38, ZN => p_14_port);
   U93 : MUX2_X1 port map( A => net29998, B => n50, S => A(15), Z => n41);
   U94 : MUX2_X1 port map( A => n88, B => net30001, S => A(14), Z => n40);
   U95 : NAND3_X1 port map( A1 => n41, A2 => n72, A3 => n40, ZN => p_15_port);
   U96 : MUX2_X1 port map( A => n58, B => n70, S => A(16), Z => n43);
   U97 : MUX2_X1 port map( A => n88, B => net30001, S => A(15), Z => n42);
   U98 : NAND3_X1 port map( A1 => n43, A2 => n72, A3 => n42, ZN => p_16_port);
   U99 : MUX2_X1 port map( A => n58, B => n9, S => A(17), Z => n45);
   U100 : MUX2_X1 port map( A => n88, B => net30001, S => A(16), Z => n44);
   U101 : NAND3_X1 port map( A1 => n45, A2 => net42472, A3 => n44, ZN => 
                           p_17_port);
   U102 : MUX2_X1 port map( A => n88, B => net30001, S => A(17), Z => n47);
   U103 : NAND2_X1 port map( A1 => n8, A2 => net30033, ZN => n50);
   U104 : MUX2_X1 port map( A => net29998, B => n50, S => A(18), Z => n46);
   U105 : NAND3_X1 port map( A1 => n47, A2 => net42472, A3 => n46, ZN => 
                           p_18_port);
   U106 : MUX2_X1 port map( A => n88, B => net30001, S => A(18), Z => n49);
   U107 : MUX2_X1 port map( A => net29998, B => n50, S => A(19), Z => n48);
   U108 : NAND3_X1 port map( A1 => n49, A2 => n72, A3 => n48, ZN => p_19_port);
   U109 : MUX2_X1 port map( A => net29998, B => n50, S => A(20), Z => n52);
   U110 : MUX2_X1 port map( A => n88, B => net30001, S => A(19), Z => n51);
   U112 : MUX2_X1 port map( A => net29998, B => n50, S => A(22), Z => n53);
   U113 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => p_22_port);
   U114 : MUX2_X1 port map( A => net29998, B => net30010, S => A(23), Z => n55)
                           ;
   U115 : NAND3_X1 port map( A1 => n55, A2 => net30022, A3 => net42472, ZN => 
                           p_23_port);
   U116 : MUX2_X1 port map( A => n88, B => net30001, S => A(23), Z => n57);
   U118 : NAND3_X1 port map( A1 => n57, A2 => n72, A3 => net29998, ZN => 
                           p_24_port);
   U121 : NAND3_X1 port map( A1 => n88, A2 => net42472, A3 => n58, ZN => 
                           p_25_port);
   U127 : NAND3_X1 port map( A1 => net29998, A2 => n72, A3 => n88, ZN => 
                           p_27_port);
   U133 : NAND3_X1 port map( A1 => n58, A2 => n72, A3 => n88, ZN => p_29_port);
   U136 : NAND3_X1 port map( A1 => n88, A2 => net42472, A3 => n58, ZN => 
                           p_30_port);
   U139 : NAND3_X1 port map( A1 => n88, A2 => n72, A3 => n58, ZN => p_31_port);
   U11 : INV_X1 port map( A => net34028, ZN => n58);
   U4 : NAND3_X1 port map( A1 => n52, A2 => n51, A3 => n72, ZN => p_20_port);
   U6 : NAND2_X1 port map( A1 => net29998, A2 => n87, ZN => p_26_port);
   U20 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n83);
   U22 : AND3_X1 port map( A1 => b(2), A2 => n78, A3 => n1, ZN => net33339);
   U27 : OAI21_X1 port map( B1 => net33339, B2 => A(20), A => n86, ZN => 
                           net30030);
   U28 : NAND2_X1 port map( A1 => net30001, A2 => A(20), ZN => n86);
   U30 : NAND2_X1 port map( A1 => n58, A2 => n88, ZN => p_32_port);
   U32 : MUX2_X1 port map( A => n88, B => net30001, S => A(22), Z => net30022);
   U33 : MUX2_X1 port map( A => n88, B => net30001, S => A(2), Z => n17);
   U43 : MUX2_X1 port map( A => n88, B => net30001, S => A(13), Z => n38);
   U57 : AND2_X1 port map( A1 => n72, A2 => n88, ZN => n87);
   U26 : INV_X1 port map( A => b(1), ZN => n78);
   U9 : AND2_X1 port map( A1 => net30075, A2 => b(2), ZN => net34028);
   U19 : NAND2_X1 port map( A1 => net34028, A2 => net30077, ZN => net42472);
   U3 : NAND2_X2 port map( A1 => b(0), A2 => b(1), ZN => net30001);
   U5 : NAND2_X1 port map( A1 => b(2), A2 => n83, ZN => net29998);
   U7 : NAND2_X2 port map( A1 => net34028, A2 => net30077, ZN => n72);
   U10 : INV_X2 port map( A => net33339, ZN => n88);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_14 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_14;

architecture SYN_beh of ENC_14 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n6, n14, n15, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, 
      n65, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n84, n86, n93, n96, n99, n101, n105, n113 : std_logic;

begin
   
   U9 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n31);
   U10 : NAND2_X1 port map( A1 => b(0), A2 => n113, ZN => n2);
   U11 : NAND2_X1 port map( A1 => n29, A2 => b(1), ZN => n3);
   U12 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => n71);
   U21 : NAND2_X1 port map( A1 => n27, A2 => n76, ZN => n6);
   U32 : AND2_X1 port map( A1 => n31, A2 => b(2), ZN => n15);
   U33 : NAND2_X1 port map( A1 => n14, A2 => n113, ZN => n96);
   U34 : INV_X1 port map( A => b(2), ZN => n76);
   U36 : INV_X1 port map( A => b(0), ZN => n29);
   U39 : NAND2_X1 port map( A1 => b(2), A2 => n84, ZN => n30);
   U41 : MUX2_X1 port map( A => n30, B => n99, S => A(0), Z => n28);
   U42 : OAI211_X1 port map( C1 => n76, C2 => n84, A => n96, B => n28, ZN => 
                           p(0));
   U43 : MUX2_X1 port map( A => n96, B => n84, S => A(0), Z => n33);
   U46 : MUX2_X1 port map( A => n105, B => n99, S => A(1), Z => n32);
   U47 : NAND3_X1 port map( A1 => n33, A2 => n101, A3 => n32, ZN => p(1));
   U48 : MUX2_X1 port map( A => n96, B => n84, S => A(1), Z => n35);
   U49 : MUX2_X1 port map( A => n105, B => n99, S => A(2), Z => n34);
   U50 : NAND3_X1 port map( A1 => n35, A2 => n101, A3 => n34, ZN => p(2));
   U51 : MUX2_X1 port map( A => n93, B => n84, S => A(2), Z => n37);
   U52 : MUX2_X1 port map( A => n105, B => n6, S => A(3), Z => n36);
   U53 : NAND3_X1 port map( A1 => n37, A2 => n101, A3 => n36, ZN => p(3));
   U54 : MUX2_X1 port map( A => n93, B => n84, S => A(3), Z => n39);
   U55 : MUX2_X1 port map( A => n105, B => n99, S => A(4), Z => n38);
   U56 : NAND3_X1 port map( A1 => n39, A2 => n101, A3 => n38, ZN => p(4));
   U57 : MUX2_X1 port map( A => n93, B => n84, S => A(4), Z => n41);
   U58 : MUX2_X1 port map( A => n105, B => n99, S => A(5), Z => n40);
   U59 : NAND3_X1 port map( A1 => n41, A2 => n101, A3 => n40, ZN => p(5));
   U60 : MUX2_X1 port map( A => n93, B => n84, S => A(5), Z => n43);
   U61 : MUX2_X1 port map( A => n105, B => n6, S => A(6), Z => n42);
   U62 : NAND3_X1 port map( A1 => n43, A2 => n101, A3 => n42, ZN => p(6));
   U63 : MUX2_X1 port map( A => n93, B => n84, S => A(6), Z => n45);
   U64 : MUX2_X1 port map( A => n105, B => n99, S => A(7), Z => n44);
   U65 : NAND3_X1 port map( A1 => n45, A2 => n101, A3 => n44, ZN => p(7));
   U66 : MUX2_X1 port map( A => n96, B => n84, S => A(7), Z => n47);
   U67 : MUX2_X1 port map( A => n105, B => n99, S => A(8), Z => n46);
   U68 : NAND3_X1 port map( A1 => n46, A2 => n101, A3 => n47, ZN => p(8));
   U69 : MUX2_X1 port map( A => n93, B => n84, S => A(8), Z => n49);
   U70 : MUX2_X1 port map( A => n105, B => n99, S => A(9), Z => n48);
   U71 : NAND3_X1 port map( A1 => n49, A2 => n101, A3 => n48, ZN => p(9));
   U72 : MUX2_X1 port map( A => n96, B => n84, S => A(9), Z => n51);
   U73 : MUX2_X1 port map( A => n105, B => n6, S => A(10), Z => n50);
   U74 : NAND3_X1 port map( A1 => n51, A2 => n101, A3 => n50, ZN => p(10));
   U75 : MUX2_X1 port map( A => n93, B => n84, S => A(10), Z => n53);
   U76 : MUX2_X1 port map( A => n105, B => n99, S => A(11), Z => n52);
   U77 : NAND3_X1 port map( A1 => n53, A2 => n101, A3 => n52, ZN => p(11));
   U78 : MUX2_X1 port map( A => n93, B => n84, S => A(11), Z => n55);
   U79 : MUX2_X1 port map( A => n105, B => n99, S => A(12), Z => n54);
   U80 : NAND3_X1 port map( A1 => n55, A2 => n101, A3 => n54, ZN => p(12));
   U81 : MUX2_X1 port map( A => n96, B => n84, S => A(12), Z => n57);
   U82 : MUX2_X1 port map( A => n105, B => n99, S => A(13), Z => n56);
   U83 : NAND3_X1 port map( A1 => n57, A2 => n101, A3 => n56, ZN => p(13));
   U84 : MUX2_X1 port map( A => n93, B => n84, S => A(13), Z => n59);
   U85 : MUX2_X1 port map( A => n105, B => n99, S => A(14), Z => n58);
   U86 : NAND3_X1 port map( A1 => n59, A2 => n101, A3 => n58, ZN => p(14));
   U87 : MUX2_X1 port map( A => n96, B => n84, S => A(14), Z => n61);
   U88 : MUX2_X1 port map( A => n105, B => n99, S => A(15), Z => n60);
   U89 : NAND3_X1 port map( A1 => n61, A2 => n101, A3 => n60, ZN => p(15));
   U90 : MUX2_X1 port map( A => n86, B => n84, S => A(15), Z => n63);
   U91 : MUX2_X1 port map( A => n105, B => n6, S => A(16), Z => n62);
   U92 : NAND3_X1 port map( A1 => n63, A2 => n101, A3 => n62, ZN => p(16));
   U93 : MUX2_X1 port map( A => n105, B => n99, S => A(17), Z => n65);
   U94 : MUX2_X1 port map( A => n96, B => n84, S => A(16), Z => n64);
   U95 : NAND3_X1 port map( A1 => n65, A2 => n101, A3 => n64, ZN => p(17));
   U96 : MUX2_X1 port map( A => n93, B => n84, S => A(17), Z => n68);
   U97 : MUX2_X1 port map( A => n105, B => n99, S => A(18), Z => n67);
   U98 : NAND3_X1 port map( A1 => n68, A2 => n101, A3 => n67, ZN => p(18));
   U99 : MUX2_X1 port map( A => n105, B => n99, S => A(19), Z => n70);
   U100 : MUX2_X1 port map( A => n93, B => n84, S => A(18), Z => n69);
   U101 : NAND3_X1 port map( A1 => n70, A2 => n101, A3 => n69, ZN => p(19));
   U102 : MUX2_X1 port map( A => n86, B => n84, S => A(19), Z => n73);
   U103 : NAND2_X1 port map( A1 => n71, A2 => n76, ZN => n81);
   U104 : MUX2_X1 port map( A => n105, B => n81, S => A(20), Z => n72);
   U105 : NAND3_X1 port map( A1 => n72, A2 => n101, A3 => n73, ZN => p(20));
   U106 : MUX2_X1 port map( A => n86, B => n84, S => A(20), Z => n75);
   U107 : MUX2_X1 port map( A => n105, B => n6, S => A(21), Z => n74);
   U108 : NAND3_X1 port map( A1 => n75, A2 => n101, A3 => n74, ZN => p(21));
   U109 : MUX2_X1 port map( A => n105, B => n81, S => A(22), Z => n78);
   U110 : MUX2_X1 port map( A => n86, B => n84, S => A(21), Z => n77);
   U112 : MUX2_X1 port map( A => n105, B => n81, S => A(23), Z => n80);
   U113 : MUX2_X1 port map( A => n96, B => n84, S => A(22), Z => n79);
   U114 : NAND3_X1 port map( A1 => n80, A2 => n79, A3 => n101, ZN => p(23));
   U116 : MUX2_X1 port map( A => n86, B => n84, S => A(23), Z => n82);
   U117 : NAND3_X1 port map( A1 => n82, A2 => n101, A3 => n105, ZN => p(24));
   U120 : NAND3_X1 port map( A1 => n93, A2 => n101, A3 => n105, ZN => p(25));
   U123 : NAND3_X1 port map( A1 => n93, A2 => n105, A3 => n101, ZN => p(26));
   U126 : NAND3_X1 port map( A1 => n105, A2 => n101, A3 => n93, ZN => p(27));
   U129 : NAND3_X1 port map( A1 => n96, A2 => n105, A3 => n101, ZN => p(28));
   U132 : NAND3_X1 port map( A1 => n93, A2 => n101, A3 => n105, ZN => p(29));
   U135 : NAND3_X1 port map( A1 => n93, A2 => n101, A3 => n105, ZN => p(30));
   U138 : NAND3_X1 port map( A1 => n96, A2 => n101, A3 => n105, ZN => p(31));
   U140 : NAND2_X1 port map( A1 => n105, A2 => n96, ZN => p(32));
   U14 : XNOR2_X1 port map( A => b(0), B => n113, ZN => n27);
   U15 : NAND2_X1 port map( A1 => n14, A2 => n113, ZN => n86);
   U17 : NAND3_X1 port map( A1 => n77, A2 => n78, A3 => n101, ZN => p(22));
   U7 : AND2_X1 port map( A1 => n29, A2 => b(2), ZN => n14);
   U13 : NAND2_X1 port map( A1 => n76, A2 => n27, ZN => n99);
   U16 : INV_X1 port map( A => b(1), ZN => n113);
   U3 : NAND2_X2 port map( A1 => b(0), A2 => b(1), ZN => n84);
   U4 : NAND2_X2 port map( A1 => n31, A2 => b(2), ZN => n105);
   U5 : NAND2_X2 port map( A1 => n15, A2 => n30, ZN => n101);
   U6 : NAND2_X2 port map( A1 => n14, A2 => n113, ZN => n93);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_15 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_15;

architecture SYN_beh of ENC_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n5, n6, n9, n11, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, 
      n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60
      , n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, 
      n75, n76, n79, n83, n85, n90, n94, n98, n101, n105, n109, n110, n112, 
      n114, n115, n118, n119 : std_logic;

begin
   
   U9 : NAND2_X1 port map( A1 => n75, A2 => n114, ZN => n5);
   U10 : NAND2_X1 port map( A1 => n83, A2 => A(23), ZN => n6);
   U11 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => n72);
   U15 : NAND2_X1 port map( A1 => n11, A2 => n105, ZN => n76);
   U19 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => n9);
   U31 : NAND2_X1 port map( A1 => b(2), A2 => n98, ZN => n23);
   U34 : MUX2_X1 port map( A => n23, B => n1, S => A(0), Z => n22);
   U35 : OAI211_X1 port map( C1 => n61, C2 => n85, A => n110, B => n22, ZN => 
                           p(0));
   U37 : MUX2_X1 port map( A => n109, B => n98, S => A(0), Z => n26);
   U39 : MUX2_X1 port map( A => n75, B => n1, S => A(1), Z => n25);
   U40 : NAND3_X1 port map( A1 => n26, A2 => n118, A3 => n25, ZN => p(1));
   U41 : MUX2_X1 port map( A => n109, B => n98, S => A(1), Z => n28);
   U42 : MUX2_X1 port map( A => n75, B => n1, S => A(2), Z => n27);
   U43 : NAND3_X1 port map( A1 => n28, A2 => n118, A3 => n27, ZN => p(2));
   U44 : MUX2_X1 port map( A => n76, B => n85, S => A(2), Z => n30);
   U45 : MUX2_X1 port map( A => n101, B => n1, S => A(3), Z => n29);
   U46 : NAND3_X1 port map( A1 => n30, A2 => n118, A3 => n29, ZN => p(3));
   U47 : MUX2_X1 port map( A => n110, B => n85, S => A(3), Z => n32);
   U48 : MUX2_X1 port map( A => n101, B => n1, S => A(4), Z => n31);
   U49 : NAND3_X1 port map( A1 => n32, A2 => n118, A3 => n31, ZN => p(4));
   U50 : MUX2_X1 port map( A => n76, B => n85, S => A(4), Z => n34);
   U51 : MUX2_X1 port map( A => n75, B => n1, S => A(5), Z => n33);
   U52 : NAND3_X1 port map( A1 => n34, A2 => n118, A3 => n33, ZN => p(5));
   U53 : MUX2_X1 port map( A => n109, B => n98, S => A(5), Z => n36);
   U54 : MUX2_X1 port map( A => n101, B => n1, S => A(6), Z => n35);
   U55 : NAND3_X1 port map( A1 => n36, A2 => n118, A3 => n35, ZN => p(6));
   U56 : MUX2_X1 port map( A => n76, B => n85, S => A(6), Z => n38);
   U57 : MUX2_X1 port map( A => n101, B => n1, S => A(7), Z => n37);
   U58 : NAND3_X1 port map( A1 => n38, A2 => n118, A3 => n37, ZN => p(7));
   U59 : MUX2_X1 port map( A => n109, B => n98, S => A(7), Z => n40);
   U60 : MUX2_X1 port map( A => n101, B => n94, S => A(8), Z => n39);
   U61 : NAND3_X1 port map( A1 => n40, A2 => n118, A3 => n39, ZN => p(8));
   U62 : MUX2_X1 port map( A => n110, B => n98, S => A(8), Z => n42);
   U63 : MUX2_X1 port map( A => n101, B => n94, S => A(9), Z => n41);
   U64 : NAND3_X1 port map( A1 => n42, A2 => n118, A3 => n41, ZN => p(9));
   U65 : MUX2_X1 port map( A => n76, B => n98, S => A(9), Z => n44);
   U66 : MUX2_X1 port map( A => n101, B => n1, S => A(10), Z => n43);
   U67 : NAND3_X1 port map( A1 => n44, A2 => n118, A3 => n43, ZN => p(10));
   U68 : MUX2_X1 port map( A => n76, B => n98, S => A(10), Z => n46);
   U69 : MUX2_X1 port map( A => n101, B => n1, S => A(11), Z => n45);
   U70 : NAND3_X1 port map( A1 => n46, A2 => n118, A3 => n45, ZN => p(11));
   U71 : MUX2_X1 port map( A => n109, B => n98, S => A(11), Z => n48);
   U72 : MUX2_X1 port map( A => n101, B => n1, S => A(12), Z => n47);
   U73 : NAND3_X1 port map( A1 => n48, A2 => n118, A3 => n47, ZN => p(12));
   U74 : MUX2_X1 port map( A => n110, B => n85, S => A(12), Z => n50);
   U75 : MUX2_X1 port map( A => n101, B => n1, S => A(13), Z => n49);
   U76 : NAND3_X1 port map( A1 => n50, A2 => n118, A3 => n49, ZN => p(13));
   U77 : MUX2_X1 port map( A => n76, B => n98, S => A(13), Z => n52);
   U78 : MUX2_X1 port map( A => n101, B => n94, S => A(14), Z => n51);
   U79 : NAND3_X1 port map( A1 => n52, A2 => n118, A3 => n51, ZN => p(14));
   U80 : MUX2_X1 port map( A => n110, B => n98, S => A(14), Z => n54);
   U81 : MUX2_X1 port map( A => n101, B => n1, S => A(15), Z => n53);
   U82 : NAND3_X1 port map( A1 => n54, A2 => n118, A3 => n53, ZN => p(15));
   U83 : MUX2_X1 port map( A => n76, B => n98, S => A(15), Z => n56);
   U84 : MUX2_X1 port map( A => n101, B => n1, S => A(16), Z => n55);
   U85 : NAND3_X1 port map( A1 => n55, A2 => n118, A3 => n56, ZN => p(16));
   U86 : MUX2_X1 port map( A => n110, B => n98, S => A(16), Z => n58);
   U87 : MUX2_X1 port map( A => n101, B => n94, S => A(17), Z => n57);
   U88 : NAND3_X1 port map( A1 => n58, A2 => n118, A3 => n57, ZN => p(17));
   U89 : MUX2_X1 port map( A => n90, B => n98, S => A(17), Z => n60);
   U90 : MUX2_X1 port map( A => n101, B => n1, S => A(18), Z => n59);
   U91 : NAND3_X1 port map( A1 => n60, A2 => n118, A3 => n59, ZN => p(18));
   U92 : MUX2_X1 port map( A => n109, B => n98, S => A(18), Z => n64);
   U93 : XOR2_X1 port map( A => b(0), B => b(1), Z => n62);
   U94 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => n83);
   U95 : MUX2_X1 port map( A => n101, B => n9, S => A(19), Z => n63);
   U96 : NAND3_X1 port map( A1 => n64, A2 => n118, A3 => n63, ZN => p(19));
   U97 : MUX2_X1 port map( A => n76, B => n98, S => A(19), Z => n66);
   U98 : MUX2_X1 port map( A => n101, B => n1, S => A(20), Z => n65);
   U99 : NAND3_X1 port map( A1 => n66, A2 => n118, A3 => n65, ZN => p(20));
   U100 : MUX2_X1 port map( A => n110, B => n98, S => A(20), Z => n68);
   U101 : MUX2_X1 port map( A => n101, B => n1, S => A(21), Z => n67);
   U102 : NAND3_X1 port map( A1 => n68, A2 => n118, A3 => n67, ZN => p(21));
   U103 : MUX2_X1 port map( A => n110, B => n98, S => A(21), Z => n71);
   U104 : NAND2_X1 port map( A1 => b(2), A2 => n69, ZN => n75);
   U105 : MUX2_X1 port map( A => n75, B => n9, S => A(22), Z => n70);
   U106 : NAND3_X1 port map( A1 => n71, A2 => n70, A3 => n118, ZN => p(22));
   U107 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n85);
   U108 : MUX2_X1 port map( A => n79, B => n85, S => A(22), Z => n73);
   U109 : NAND3_X1 port map( A1 => n72, A2 => n73, A3 => n118, ZN => p(23));
   U115 : NAND3_X1 port map( A1 => n75, A2 => n118, A3 => n90, ZN => p(25));
   U117 : NAND2_X1 port map( A1 => n11, A2 => n105, ZN => n79);
   U119 : NAND3_X1 port map( A1 => n75, A2 => n118, A3 => n109, ZN => p(26));
   U122 : NAND3_X1 port map( A1 => n109, A2 => n118, A3 => n75, ZN => p(27));
   U125 : NAND3_X1 port map( A1 => n75, A2 => n90, A3 => n118, ZN => p(28));
   U128 : NAND3_X1 port map( A1 => n90, A2 => n118, A3 => n101, ZN => p(29));
   U136 : NAND2_X1 port map( A1 => n101, A2 => n90, ZN => p(32));
   U3 : XNOR2_X1 port map( A => n105, B => b(0), ZN => n21);
   U12 : NAND2_X1 port map( A1 => n11, A2 => n105, ZN => n90);
   U16 : NAND2_X1 port map( A1 => n11, A2 => n105, ZN => n109);
   U17 : NAND2_X1 port map( A1 => n11, A2 => n105, ZN => n110);
   U21 : NAND2_X1 port map( A1 => n98, A2 => A(23), ZN => n112);
   U22 : INV_X1 port map( A => b(0), ZN => n115);
   U26 : INV_X1 port map( A => A(23), ZN => n114);
   U27 : NAND3_X1 port map( A1 => n74, A2 => n118, A3 => n75, ZN => p(24));
   U30 : AND2_X1 port map( A1 => n115, A2 => b(2), ZN => n11);
   U13 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n98);
   U131 : NAND3_X1 port map( A1 => n90, A2 => n118, A3 => n101, ZN => p(30));
   U134 : NAND3_X1 port map( A1 => n90, A2 => n118, A3 => n101, ZN => p(31));
   U4 : NAND2_X1 port map( A1 => n21, A2 => n61, ZN => n1);
   U5 : NAND2_X1 port map( A1 => b(2), A2 => n69, ZN => n101);
   U6 : NAND3_X2 port map( A1 => b(0), A2 => b(2), A3 => b(1), ZN => n118);
   U7 : OR2_X1 port map( A1 => b(0), A2 => b(1), ZN => n69);
   U8 : INV_X1 port map( A => b(1), ZN => n105);
   U18 : INV_X1 port map( A => b(2), ZN => n61);
   U20 : NAND2_X1 port map( A1 => n21, A2 => n61, ZN => n94);
   U23 : NAND2_X1 port map( A1 => n119, A2 => n112, ZN => n74);
   U24 : NAND2_X1 port map( A1 => n114, A2 => n79, ZN => n119);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_16 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_16;

architecture SYN_beh of ENC_16 is

   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal p_32_port, p_31_port, p_29_port, p_28_port, p_27_port, p_26_port, 
      p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, p_20_port, 
      p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, p_14_port, 
      p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port, p_7_port,
      p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, p_0_port, n7,
      n10, n11, n12, n13, n27, n28, n29, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
      n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n86, n88, n98, n100, n102, n108 : std_logic;

begin
   p <= ( p_32_port, p_31_port, p_31_port, p_29_port, p_28_port, p_27_port, 
      p_26_port, p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, 
      p_20_port, p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, 
      p_14_port, p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port
      , p_7_port, p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, 
      p_0_port );
   
   U11 : NAND2_X1 port map( A1 => n12, A2 => b(2), ZN => n88);
   U27 : XNOR2_X1 port map( A => b(0), B => n108, ZN => n11);
   U28 : NAND2_X1 port map( A1 => n7, A2 => n108, ZN => n12);
   U29 : NAND2_X1 port map( A1 => n11, A2 => n63, ZN => n13);
   U31 : NAND2_X1 port map( A1 => n11, A2 => n63, ZN => n69);
   U33 : INV_X1 port map( A => b(2), ZN => n63);
   U34 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n28);
   U38 : NAND2_X1 port map( A1 => b(2), A2 => n28, ZN => n29);
   U39 : MUX2_X1 port map( A => n29, B => n13, S => A(0), Z => n27);
   U40 : OAI211_X1 port map( C1 => n63, C2 => n10, A => n102, B => n27, ZN => 
                           p_0_port);
   U41 : MUX2_X1 port map( A => n102, B => n10, S => A(0), Z => n33);
   U43 : NAND2_X1 port map( A1 => n7, A2 => n108, ZN => n62);
   U44 : MUX2_X1 port map( A => n82, B => n13, S => A(1), Z => n32);
   U45 : NAND3_X1 port map( A1 => n33, A2 => n100, A3 => n32, ZN => p_1_port);
   U46 : MUX2_X1 port map( A => n102, B => n10, S => A(1), Z => n35);
   U47 : MUX2_X1 port map( A => n82, B => n13, S => A(2), Z => n34);
   U48 : NAND3_X1 port map( A1 => n34, A2 => n100, A3 => n35, ZN => p_2_port);
   U49 : MUX2_X1 port map( A => n102, B => n10, S => A(2), Z => n37);
   U50 : MUX2_X1 port map( A => n82, B => n69, S => A(3), Z => n36);
   U51 : NAND3_X1 port map( A1 => n37, A2 => n100, A3 => n36, ZN => p_3_port);
   U52 : MUX2_X1 port map( A => n102, B => n10, S => A(3), Z => n39);
   U53 : MUX2_X1 port map( A => n82, B => n13, S => A(4), Z => n38);
   U54 : NAND3_X1 port map( A1 => n39, A2 => n100, A3 => n38, ZN => p_4_port);
   U55 : MUX2_X1 port map( A => n102, B => n10, S => A(4), Z => n41);
   U56 : MUX2_X1 port map( A => n86, B => n69, S => A(5), Z => n40);
   U57 : NAND3_X1 port map( A1 => n41, A2 => n100, A3 => n40, ZN => p_5_port);
   U58 : MUX2_X1 port map( A => n102, B => n10, S => A(5), Z => n43);
   U59 : MUX2_X1 port map( A => n82, B => n13, S => A(6), Z => n42);
   U60 : NAND3_X1 port map( A1 => n43, A2 => n100, A3 => n42, ZN => p_6_port);
   U61 : MUX2_X1 port map( A => n102, B => n10, S => A(6), Z => n45);
   U62 : MUX2_X1 port map( A => n82, B => n69, S => A(7), Z => n44);
   U63 : NAND3_X1 port map( A1 => n45, A2 => n100, A3 => n44, ZN => p_7_port);
   U64 : MUX2_X1 port map( A => n102, B => n10, S => A(7), Z => n47);
   U65 : MUX2_X1 port map( A => n86, B => n13, S => A(8), Z => n46);
   U66 : NAND3_X1 port map( A1 => n47, A2 => n100, A3 => n46, ZN => p_8_port);
   U67 : MUX2_X1 port map( A => n102, B => n10, S => A(8), Z => n49);
   U68 : MUX2_X1 port map( A => n86, B => n69, S => A(9), Z => n48);
   U69 : NAND3_X1 port map( A1 => n49, A2 => n100, A3 => n48, ZN => p_9_port);
   U70 : MUX2_X1 port map( A => n102, B => n10, S => A(9), Z => n51);
   U71 : MUX2_X1 port map( A => n82, B => n69, S => A(10), Z => n50);
   U72 : NAND3_X1 port map( A1 => n51, A2 => n100, A3 => n50, ZN => p_10_port);
   U73 : MUX2_X1 port map( A => n82, B => n13, S => A(11), Z => n53);
   U74 : MUX2_X1 port map( A => n102, B => n10, S => A(10), Z => n52);
   U75 : NAND3_X1 port map( A1 => n53, A2 => n100, A3 => n52, ZN => p_11_port);
   U76 : MUX2_X1 port map( A => n102, B => n10, S => A(11), Z => n55);
   U77 : MUX2_X1 port map( A => n86, B => n69, S => A(12), Z => n54);
   U78 : NAND3_X1 port map( A1 => n55, A2 => n100, A3 => n54, ZN => p_12_port);
   U79 : MUX2_X1 port map( A => n86, B => n13, S => A(13), Z => n57);
   U80 : MUX2_X1 port map( A => n102, B => n10, S => A(12), Z => n56);
   U81 : NAND3_X1 port map( A1 => n100, A2 => n57, A3 => n56, ZN => p_13_port);
   U82 : MUX2_X1 port map( A => n102, B => n10, S => A(13), Z => n59);
   U83 : MUX2_X1 port map( A => n82, B => n13, S => A(14), Z => n58);
   U84 : NAND3_X1 port map( A1 => n59, A2 => n100, A3 => n58, ZN => p_14_port);
   U85 : MUX2_X1 port map( A => n86, B => n69, S => A(15), Z => n61);
   U86 : MUX2_X1 port map( A => n102, B => n10, S => A(14), Z => n60);
   U87 : NAND3_X1 port map( A1 => n61, A2 => n100, A3 => n60, ZN => p_15_port);
   U88 : NAND2_X1 port map( A1 => n12, A2 => b(2), ZN => n84);
   U89 : XOR2_X1 port map( A => b(0), B => b(1), Z => n64);
   U90 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => n98);
   U91 : MUX2_X1 port map( A => n82, B => n98, S => A(16), Z => n66);
   U92 : MUX2_X1 port map( A => n102, B => n10, S => A(15), Z => n65);
   U93 : NAND3_X1 port map( A1 => n66, A2 => n100, A3 => n65, ZN => p_16_port);
   U94 : MUX2_X1 port map( A => n82, B => n98, S => A(17), Z => n68);
   U95 : MUX2_X1 port map( A => n102, B => n10, S => A(16), Z => n67);
   U96 : NAND3_X1 port map( A1 => n68, A2 => n100, A3 => n67, ZN => p_17_port);
   U97 : MUX2_X1 port map( A => n102, B => n10, S => A(17), Z => n71);
   U98 : MUX2_X1 port map( A => n86, B => n13, S => A(18), Z => n70);
   U99 : NAND3_X1 port map( A1 => n71, A2 => n100, A3 => n70, ZN => p_18_port);
   U100 : MUX2_X1 port map( A => n88, B => n98, S => A(19), Z => n73);
   U101 : MUX2_X1 port map( A => n102, B => n10, S => A(18), Z => n72);
   U102 : NAND3_X1 port map( A1 => n73, A2 => n100, A3 => n72, ZN => p_19_port)
                           ;
   U103 : MUX2_X1 port map( A => n102, B => n10, S => A(19), Z => n75);
   U104 : MUX2_X1 port map( A => n86, B => n69, S => A(20), Z => n74);
   U105 : NAND3_X1 port map( A1 => n75, A2 => n100, A3 => n74, ZN => p_20_port)
                           ;
   U106 : MUX2_X1 port map( A => n102, B => n10, S => A(20), Z => n77);
   U107 : MUX2_X1 port map( A => n82, B => n13, S => A(21), Z => n76);
   U108 : NAND3_X1 port map( A1 => n77, A2 => n100, A3 => n76, ZN => p_21_port)
                           ;
   U109 : MUX2_X1 port map( A => n102, B => n10, S => A(21), Z => n79);
   U110 : MUX2_X1 port map( A => n84, B => n69, S => A(22), Z => n78);
   U111 : NAND3_X1 port map( A1 => n79, A2 => n100, A3 => n78, ZN => p_22_port)
                           ;
   U112 : MUX2_X1 port map( A => n102, B => n10, S => A(22), Z => n81);
   U113 : MUX2_X1 port map( A => n88, B => n69, S => A(23), Z => n80);
   U114 : NAND3_X1 port map( A1 => n81, A2 => n100, A3 => n80, ZN => p_23_port)
                           ;
   U115 : MUX2_X1 port map( A => n102, B => n10, S => A(23), Z => n83);
   U117 : NAND3_X1 port map( A1 => n83, A2 => n82, A3 => n100, ZN => p_24_port)
                           ;
   U120 : NAND3_X1 port map( A1 => n84, A2 => n102, A3 => n100, ZN => p_25_port
                           );
   U123 : NAND3_X1 port map( A1 => n102, A2 => n86, A3 => n100, ZN => p_26_port
                           );
   U128 : NAND3_X1 port map( A1 => n102, A2 => n100, A3 => n84, ZN => p_28_port
                           );
   U131 : NAND3_X1 port map( A1 => n86, A2 => n100, A3 => n102, ZN => p_29_port
                           );
   U137 : NAND3_X1 port map( A1 => n102, A2 => n100, A3 => n86, ZN => p_31_port
                           );
   U139 : NAND2_X1 port map( A1 => n86, A2 => n102, ZN => p_32_port);
   U12 : NAND3_X1 port map( A1 => n100, A2 => n102, A3 => n88, ZN => p_27_port)
                           ;
   U5 : NAND2_X1 port map( A1 => n62, A2 => b(2), ZN => n86);
   U6 : NAND2_X1 port map( A1 => n62, A2 => b(2), ZN => n82);
   U3 : NAND2_X1 port map( A1 => b(0), A2 => b(1), ZN => n10);
   U10 : INV_X1 port map( A => b(0), ZN => n7);
   U14 : INV_X1 port map( A => b(1), ZN => n108);
   U4 : NAND3_X4 port map( A1 => b(2), A2 => n108, A3 => n7, ZN => n102);
   U7 : NAND2_X2 port map( A1 => n29, A2 => b(2), ZN => n100);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity ENC_0 is

   port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
         downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
         std_logic);

end ENC_0;

architecture SYN_beh of ENC_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal p_32_port, p_31_port, p_29_port, p_27_port, p_25_port, p_24_port, 
      p_23_port, p_22_port, p_21_port, p_20_port, p_19_port, p_18_port, 
      p_17_port, p_16_port, p_15_port, p_14_port, p_13_port, p_12_port, 
      p_11_port, p_10_port, p_9_port, p_8_port, p_7_port, p_6_port, p_5_port, 
      p_4_port, p_3_port, p_2_port, p_1_port, p_0_port, n7, n8, n19, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37
      , n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, 
      n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66
      , n67, n68, n70, n73, n75, n80, n84, p_30_port, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n119, n120, n122, n127 : std_logic;

begin
   p <= ( p_32_port, p_31_port, p_30_port, p_29_port, p_29_port, p_27_port, 
      p_32_port, p_25_port, p_24_port, p_23_port, p_22_port, p_21_port, 
      p_20_port, p_19_port, p_18_port, p_17_port, p_16_port, p_15_port, 
      p_14_port, p_13_port, p_12_port, p_11_port, p_10_port, p_9_port, p_8_port
      , p_7_port, p_6_port, p_5_port, p_4_port, p_3_port, p_2_port, p_1_port, 
      p_0_port );
   
   U4 : INV_X1 port map( A => b(2), ZN => n51);
   U18 : NAND2_X1 port map( A1 => b(1), A2 => n51, ZN => n7);
   U19 : NAND2_X1 port map( A1 => b(1), A2 => n51, ZN => n8);
   U23 : NAND2_X1 port map( A1 => n95, A2 => b(2), ZN => n75);
   U25 : NAND2_X1 port map( A1 => b(1), A2 => n51, ZN => n64);
   U26 : MUX2_X1 port map( A => n51, B => n7, S => A(0), Z => n19);
   U31 : MUX2_X1 port map( A => n80, B => n64, S => A(1), Z => n21);
   U34 : MUX2_X1 port map( A => n80, B => n8, S => A(2), Z => n23);
   U37 : MUX2_X1 port map( A => n80, B => n84, S => A(3), Z => n25);
   U40 : MUX2_X1 port map( A => n127, B => n7, S => A(4), Z => n27);
   U43 : MUX2_X1 port map( A => n80, B => n64, S => A(5), Z => n29);
   U46 : MUX2_X1 port map( A => n80, B => n8, S => A(6), Z => n31);
   U49 : MUX2_X1 port map( A => n127, B => n84, S => A(7), Z => n33);
   U52 : MUX2_X1 port map( A => n80, B => n8, S => A(8), Z => n35);
   U55 : MUX2_X1 port map( A => n127, B => n64, S => A(9), Z => n37);
   U58 : MUX2_X1 port map( A => n80, B => n7, S => A(10), Z => n39);
   U61 : MUX2_X1 port map( A => n80, B => n7, S => A(11), Z => n41);
   U64 : MUX2_X1 port map( A => n80, B => n8, S => A(12), Z => n43);
   U67 : MUX2_X1 port map( A => n127, B => n84, S => A(13), Z => n45);
   U70 : MUX2_X1 port map( A => n80, B => n84, S => A(14), Z => n47);
   U72 : MUX2_X1 port map( A => n80, B => n64, S => A(15), Z => n50);
   U76 : NAND2_X1 port map( A1 => b(1), A2 => n51, ZN => n84);
   U77 : MUX2_X1 port map( A => n80, B => n84, S => A(16), Z => n52);
   U80 : MUX2_X1 port map( A => n80, B => n7, S => A(17), Z => n54);
   U83 : MUX2_X1 port map( A => n80, B => n64, S => A(18), Z => n56);
   U86 : MUX2_X1 port map( A => n80, B => n8, S => A(19), Z => n58);
   U89 : MUX2_X1 port map( A => n80, B => n8, S => A(20), Z => n60);
   U92 : MUX2_X1 port map( A => n80, B => n64, S => A(21), Z => n62);
   U95 : MUX2_X1 port map( A => n80, B => n7, S => A(22), Z => n65);
   U97 : MUX2_X1 port map( A => n127, B => n64, S => A(23), Z => n68);
   U107 : NAND2_X1 port map( A1 => n95, A2 => b(2), ZN => n73);
   U126 : NAND2_X1 port map( A1 => n127, A2 => n73, ZN => p_32_port);
   U3 : NAND2_X1 port map( A1 => n63, A2 => n62, ZN => p_21_port);
   U5 : NAND2_X1 port map( A1 => n68, A2 => n67, ZN => p_23_port);
   U6 : NAND2_X1 port map( A1 => n57, A2 => n56, ZN => p_18_port);
   U7 : NAND2_X1 port map( A1 => n75, A2 => n80, ZN => p_25_port);
   U8 : NAND2_X1 port map( A1 => n70, A2 => n80, ZN => p_24_port);
   U9 : NAND2_X1 port map( A1 => n105, A2 => n107, ZN => n70);
   U10 : NAND2_X1 port map( A1 => n75, A2 => n127, ZN => p_27_port);
   U12 : NAND2_X1 port map( A1 => n42, A2 => n41, ZN => p_11_port);
   U13 : NAND2_X1 port map( A1 => n44, A2 => n43, ZN => p_12_port);
   U14 : NAND2_X1 port map( A1 => n55, A2 => n54, ZN => p_17_port);
   U15 : NAND2_X1 port map( A1 => n46, A2 => n45, ZN => p_13_port);
   U17 : NAND2_X1 port map( A1 => n53, A2 => n52, ZN => p_16_port);
   U20 : NAND2_X1 port map( A1 => n59, A2 => n58, ZN => p_19_port);
   U21 : NAND2_X1 port map( A1 => n127, A2 => n73, ZN => p_31_port);
   U24 : NAND2_X1 port map( A1 => n61, A2 => n60, ZN => p_20_port);
   U28 : NAND2_X1 port map( A1 => n75, A2 => n127, ZN => p_30_port);
   U29 : NAND2_X1 port map( A1 => n66, A2 => n65, ZN => p_22_port);
   U30 : NAND2_X1 port map( A1 => n73, A2 => n127, ZN => p_29_port);
   U32 : NAND2_X1 port map( A1 => n105, A2 => n96, ZN => n48);
   U33 : INV_X1 port map( A => A(13), ZN => n96);
   U35 : NAND2_X1 port map( A1 => n105, A2 => n97, ZN => n49);
   U36 : INV_X1 port map( A => A(14), ZN => n97);
   U38 : NAND2_X1 port map( A1 => n105, A2 => n98, ZN => n53);
   U39 : INV_X1 port map( A => A(15), ZN => n98);
   U41 : NAND2_X1 port map( A1 => n105, A2 => n99, ZN => n55);
   U42 : INV_X1 port map( A => A(16), ZN => n99);
   U44 : NAND2_X1 port map( A1 => n105, A2 => n100, ZN => n57);
   U45 : INV_X1 port map( A => A(17), ZN => n100);
   U47 : NAND2_X1 port map( A1 => n105, A2 => n101, ZN => n59);
   U48 : INV_X1 port map( A => A(18), ZN => n101);
   U50 : NAND2_X1 port map( A1 => n105, A2 => n102, ZN => n61);
   U51 : INV_X1 port map( A => A(19), ZN => n102);
   U53 : NAND2_X1 port map( A1 => n105, A2 => n103, ZN => n63);
   U54 : INV_X1 port map( A => A(20), ZN => n103);
   U56 : NAND2_X1 port map( A1 => n105, A2 => n104, ZN => n66);
   U57 : INV_X1 port map( A => A(21), ZN => n104);
   U59 : NAND2_X1 port map( A1 => n105, A2 => n106, ZN => n67);
   U60 : INV_X1 port map( A => A(22), ZN => n106);
   U63 : INV_X1 port map( A => A(23), ZN => n107);
   U65 : NAND2_X1 port map( A1 => n22, A2 => n21, ZN => p_1_port);
   U66 : NAND2_X1 port map( A1 => n48, A2 => n47, ZN => p_14_port);
   U68 : NAND2_X1 port map( A1 => n40, A2 => n39, ZN => p_10_port);
   U69 : NAND2_X1 port map( A1 => n38, A2 => n37, ZN => p_9_port);
   U71 : NAND2_X1 port map( A1 => n36, A2 => n35, ZN => p_8_port);
   U73 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => p_7_port);
   U74 : NAND2_X1 port map( A1 => n32, A2 => n31, ZN => p_6_port);
   U75 : NAND2_X1 port map( A1 => n30, A2 => n29, ZN => p_5_port);
   U78 : NAND2_X1 port map( A1 => n28, A2 => n27, ZN => p_4_port);
   U79 : NAND2_X1 port map( A1 => n26, A2 => n25, ZN => p_3_port);
   U81 : NAND2_X1 port map( A1 => n24, A2 => n23, ZN => p_2_port);
   U82 : NAND2_X1 port map( A1 => n50, A2 => n49, ZN => p_15_port);
   U84 : NAND2_X1 port map( A1 => n75, A2 => n19, ZN => p_0_port);
   U85 : NAND2_X1 port map( A1 => n105, A2 => n108, ZN => n22);
   U87 : INV_X1 port map( A => A(0), ZN => n108);
   U88 : NAND2_X1 port map( A1 => n105, A2 => n109, ZN => n24);
   U90 : INV_X1 port map( A => A(1), ZN => n109);
   U91 : NAND2_X1 port map( A1 => n105, A2 => n110, ZN => n26);
   U93 : INV_X1 port map( A => A(2), ZN => n110);
   U94 : NAND2_X1 port map( A1 => n105, A2 => n111, ZN => n28);
   U96 : INV_X1 port map( A => A(3), ZN => n111);
   U98 : NAND2_X1 port map( A1 => n105, A2 => n112, ZN => n30);
   U99 : INV_X1 port map( A => A(4), ZN => n112);
   U100 : NAND2_X1 port map( A1 => n105, A2 => n113, ZN => n32);
   U101 : INV_X1 port map( A => A(5), ZN => n113);
   U102 : NAND2_X1 port map( A1 => n105, A2 => n114, ZN => n34);
   U103 : INV_X1 port map( A => A(6), ZN => n114);
   U104 : NAND2_X1 port map( A1 => n105, A2 => n115, ZN => n36);
   U105 : INV_X1 port map( A => A(7), ZN => n115);
   U106 : NAND2_X1 port map( A1 => n105, A2 => n116, ZN => n38);
   U108 : INV_X1 port map( A => A(8), ZN => n116);
   U109 : NAND2_X1 port map( A1 => n105, A2 => n117, ZN => n40);
   U110 : INV_X1 port map( A => A(9), ZN => n117);
   U111 : NAND2_X1 port map( A1 => n105, A2 => n119, ZN => n42);
   U112 : INV_X1 port map( A => A(10), ZN => n119);
   U114 : NAND2_X1 port map( A1 => n105, A2 => n120, ZN => n44);
   U115 : INV_X1 port map( A => A(11), ZN => n120);
   U116 : NAND2_X1 port map( A1 => n105, A2 => n122, ZN => n46);
   U117 : INV_X1 port map( A => A(12), ZN => n122);
   U113 : INV_X1 port map( A => b(1), ZN => n95);
   U16 : NAND2_X2 port map( A1 => b(1), A2 => b(2), ZN => n80);
   U22 : INV_X1 port map( A => n75, ZN => n105);
   U27 : NAND2_X1 port map( A1 => b(2), A2 => b(1), ZN => n127);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity PackFP is

   port( SIGN : in std_logic;  EXP : in std_logic_vector (7 downto 0);  SIG : 
         in std_logic_vector (22 downto 0);  isNaN, isINF, isZ : in std_logic; 
         FP : out std_logic_vector (31 downto 0);  clk : in std_logic);

end PackFP;

architecture SYN_PackFP of PackFP is

   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal FP_30_port, FP_29_port, FP_28_port, FP_27_port, FP_26_port, 
      FP_25_port, FP_24_port, FP_23_port, FP_22_port, FP_21_port, FP_20_port, 
      FP_19_port, FP_18_port, FP_17_port, FP_16_port, FP_15_port, FP_14_port, 
      FP_13_port, FP_12_port, FP_11_port, FP_10_port, FP_9_port, FP_8_port, 
      FP_7_port, FP_6_port, FP_5_port, FP_4_port, FP_3_port, FP_2_port, 
      FP_1_port, FP_0_port, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n41, n64, n75, n76, n77, n78, n131, n136, n137, n_1866, n_1867, 
      n_1868 : std_logic;

begin
   FP <= ( SIGN, FP_30_port, FP_29_port, FP_28_port, FP_27_port, FP_26_port, 
      FP_25_port, FP_24_port, FP_23_port, FP_22_port, FP_21_port, FP_20_port, 
      FP_19_port, FP_18_port, FP_17_port, FP_16_port, FP_15_port, FP_14_port, 
      FP_13_port, FP_12_port, FP_11_port, FP_10_port, FP_9_port, FP_8_port, 
      FP_7_port, FP_6_port, FP_5_port, FP_4_port, FP_3_port, FP_2_port, 
      FP_1_port, FP_0_port );
   
   U7 : INV_X1 port map( A => isNaN, ZN => n64);
   U9 : AND2_X1 port map( A1 => SIG(0), A2 => n41, ZN => FP_0_port);
   U10 : AND2_X1 port map( A1 => SIG(1), A2 => n137, ZN => FP_1_port);
   U11 : AND2_X1 port map( A1 => SIG(2), A2 => n137, ZN => FP_2_port);
   U12 : AND2_X1 port map( A1 => n137, A2 => SIG(3), ZN => FP_3_port);
   U13 : AND2_X1 port map( A1 => n137, A2 => SIG(4), ZN => FP_4_port);
   U14 : AND2_X1 port map( A1 => n41, A2 => SIG(5), ZN => FP_5_port);
   U15 : AND2_X1 port map( A1 => n137, A2 => SIG(6), ZN => FP_6_port);
   U16 : AND2_X1 port map( A1 => n137, A2 => SIG(7), ZN => FP_7_port);
   U17 : AND2_X1 port map( A1 => n131, A2 => SIG(8), ZN => FP_8_port);
   U18 : AND2_X1 port map( A1 => n137, A2 => SIG(9), ZN => FP_9_port);
   U19 : AND2_X1 port map( A1 => n131, A2 => SIG(10), ZN => FP_10_port);
   U20 : AND2_X1 port map( A1 => n41, A2 => SIG(11), ZN => FP_11_port);
   U21 : AND2_X1 port map( A1 => SIG(12), A2 => n131, ZN => FP_12_port);
   U22 : AND2_X1 port map( A1 => n131, A2 => SIG(13), ZN => FP_13_port);
   U23 : AND2_X1 port map( A1 => n137, A2 => SIG(14), ZN => FP_14_port);
   U24 : AND2_X1 port map( A1 => SIG(15), A2 => n41, ZN => FP_15_port);
   U25 : AND2_X1 port map( A1 => n41, A2 => SIG(16), ZN => FP_16_port);
   U26 : AND2_X1 port map( A1 => n131, A2 => SIG(17), ZN => FP_17_port);
   U27 : AND2_X1 port map( A1 => n131, A2 => SIG(18), ZN => FP_18_port);
   U28 : AND2_X1 port map( A1 => n137, A2 => SIG(19), ZN => FP_19_port);
   U29 : AND2_X1 port map( A1 => n137, A2 => SIG(20), ZN => FP_20_port);
   U30 : AND2_X1 port map( A1 => n41, A2 => SIG(21), ZN => FP_21_port);
   U31 : NAND3_X1 port map( A1 => SIG(22), A2 => n3, A3 => n14, ZN => n4);
   U32 : NAND2_X1 port map( A1 => n75, A2 => n4, ZN => FP_22_port);
   U33 : AOI21_X1 port map( B1 => EXP(0), B2 => n14, A => n13, ZN => n6);
   U34 : INV_X1 port map( A => n6, ZN => FP_23_port);
   U35 : AOI21_X1 port map( B1 => EXP(1), B2 => n14, A => n13, ZN => n7);
   U36 : INV_X1 port map( A => n7, ZN => FP_24_port);
   U37 : AOI21_X1 port map( B1 => EXP(2), B2 => n14, A => n13, ZN => n8);
   U38 : INV_X1 port map( A => n8, ZN => FP_25_port);
   U39 : AOI21_X1 port map( B1 => EXP(3), B2 => n14, A => n13, ZN => n9);
   U40 : INV_X1 port map( A => n9, ZN => FP_26_port);
   U41 : AOI21_X1 port map( B1 => EXP(4), B2 => n14, A => n13, ZN => n10);
   U42 : INV_X1 port map( A => n10, ZN => FP_27_port);
   U43 : AOI21_X1 port map( B1 => EXP(5), B2 => n14, A => n13, ZN => n11);
   U44 : INV_X1 port map( A => n11, ZN => FP_28_port);
   U45 : AOI21_X1 port map( B1 => EXP(6), B2 => n14, A => n13, ZN => n12);
   U46 : INV_X1 port map( A => n12, ZN => FP_29_port);
   U47 : AOI21_X1 port map( B1 => EXP(7), B2 => n14, A => n13, ZN => n15);
   U48 : INV_X1 port map( A => n15, ZN => FP_30_port);
   MY_CLK_r_REG188_S1 : DFF_X1 port map( D => n64, CK => clk, Q => n78, QN => 
                           n_1866);
   MY_CLK_r_REG189_S2 : DFF_X1 port map( D => n78, CK => clk, Q => n77, QN => 
                           n_1867);
   MY_CLK_r_REG190_S3 : DFF_X1 port map( D => n77, CK => clk, Q => n76, QN => 
                           n_1868);
   MY_CLK_r_REG191_S4 : DFF_X1 port map( D => n76, CK => clk, Q => n75, QN => 
                           n136);
   U3 : AND3_X1 port map( A1 => n3, A2 => n14, A3 => n75, ZN => n131);
   U5 : AND3_X2 port map( A1 => n3, A2 => n14, A3 => n75, ZN => n137);
   U50 : INV_X1 port map( A => isINF, ZN => n3);
   U51 : OR2_X2 port map( A1 => isINF, A2 => n136, ZN => n13);
   U52 : AND3_X1 port map( A1 => n3, A2 => n14, A3 => n75, ZN => n41);
   U4 : INV_X2 port map( A => isZ, ZN => n14);

end SYN_PackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPnormalize_SIG_width28_1 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
         std_logic);

end FPnormalize_SIG_width28_1;

architecture SYN_FPnormalize of FPnormalize_SIG_width28_1 is

   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n6, n9, n11, n16, n25, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, 
      n91, n92, n93, n94, n95, n97, n98, n_1876, n_1877, n_1878, n_1879, n_1880
      , n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889,
      n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, 
      n_1899, n_1900 : std_logic;

begin
   
   U5 : XNOR2_X1 port map( A => n16, B => n60, ZN => EXP_out(6));
   U9 : XOR2_X1 port map( A => n54, B => n52, Z => EXP_out(0));
   U11 : NOR2_X1 port map( A1 => n92, A2 => n88, ZN => n6);
   U12 : XOR2_X1 port map( A => n55, B => n6, Z => EXP_out(1));
   U15 : XOR2_X1 port map( A => n56, B => n51, Z => EXP_out(2));
   U17 : NOR2_X1 port map( A1 => n89, A2 => n97, ZN => n9);
   U18 : XOR2_X1 port map( A => n57, B => n9, Z => EXP_out(3));
   U21 : XOR2_X1 port map( A => n98, B => n58, Z => EXP_out(4));
   U33 : MUX2_X1 port map( A => SIG_in(3), B => SIG_in(4), S => SIG_in(27), Z 
                           => SIG_out(3));
   U34 : MUX2_X1 port map( A => SIG_in(4), B => SIG_in(5), S => SIG_in(27), Z 
                           => SIG_out(4));
   U35 : MUX2_X1 port map( A => SIG_in(5), B => SIG_in(6), S => SIG_in(27), Z 
                           => SIG_out(5));
   U36 : MUX2_X1 port map( A => n62, B => n63, S => n52, Z => SIG_out(6));
   U37 : MUX2_X1 port map( A => n63, B => n64, S => n52, Z => SIG_out(7));
   U38 : MUX2_X1 port map( A => n64, B => n65, S => n52, Z => SIG_out(8));
   U39 : MUX2_X1 port map( A => n65, B => n66, S => n83, Z => SIG_out(9));
   U40 : MUX2_X1 port map( A => n66, B => n67, S => n83, Z => SIG_out(10));
   U41 : MUX2_X1 port map( A => n67, B => n68, S => n53, Z => SIG_out(11));
   U42 : MUX2_X1 port map( A => n68, B => n69, S => n52, Z => SIG_out(12));
   U43 : MUX2_X1 port map( A => n69, B => n70, S => n52, Z => SIG_out(13));
   U44 : MUX2_X1 port map( A => n70, B => n71, S => n52, Z => SIG_out(14));
   U45 : MUX2_X1 port map( A => n71, B => n72, S => n53, Z => SIG_out(15));
   U46 : MUX2_X1 port map( A => n72, B => n73, S => n53, Z => SIG_out(16));
   U47 : MUX2_X1 port map( A => n73, B => n74, S => n53, Z => SIG_out(17));
   U48 : MUX2_X1 port map( A => n74, B => n75, S => n53, Z => SIG_out(18));
   U49 : MUX2_X1 port map( A => n75, B => n76, S => n52, Z => SIG_out(19));
   U50 : MUX2_X1 port map( A => n76, B => n77, S => n52, Z => SIG_out(20));
   U51 : MUX2_X1 port map( A => n77, B => n78, S => n52, Z => SIG_out(21));
   U52 : MUX2_X1 port map( A => n78, B => n79, S => n52, Z => SIG_out(22));
   U53 : MUX2_X1 port map( A => n79, B => n80, S => n52, Z => SIG_out(23));
   U54 : MUX2_X1 port map( A => n80, B => n81, S => n53, Z => SIG_out(24));
   U55 : MUX2_X1 port map( A => n81, B => n82, S => n53, Z => SIG_out(25));
   U57 : NAND2_X1 port map( A1 => n91, A2 => n92, ZN => SIG_out(26));
   MY_CLK_r_REG205_S4 : DFF_X1 port map( D => SIG_in(27), CK => clk, Q => n83, 
                           QN => n92);
   MY_CLK_r_REG212_S4 : DFF_X1 port map( D => SIG_in(26), CK => clk, Q => n82, 
                           QN => n91);
   MY_CLK_r_REG213_S4 : DFF_X1 port map( D => SIG_in(25), CK => clk, Q => n81, 
                           QN => n_1876);
   MY_CLK_r_REG219_S4 : DFF_X1 port map( D => SIG_in(24), CK => clk, Q => n80, 
                           QN => n_1877);
   MY_CLK_r_REG214_S4 : DFF_X1 port map( D => SIG_in(23), CK => clk, Q => n79, 
                           QN => n_1878);
   MY_CLK_r_REG217_S4 : DFF_X1 port map( D => SIG_in(22), CK => clk, Q => n78, 
                           QN => n_1879);
   MY_CLK_r_REG216_S4 : DFF_X1 port map( D => SIG_in(21), CK => clk, Q => n77, 
                           QN => n_1880);
   MY_CLK_r_REG218_S4 : DFF_X1 port map( D => SIG_in(20), CK => clk, Q => n76, 
                           QN => n_1881);
   MY_CLK_r_REG215_S4 : DFF_X1 port map( D => SIG_in(19), CK => clk, Q => n75, 
                           QN => n_1882);
   MY_CLK_r_REG220_S4 : DFF_X1 port map( D => SIG_in(18), CK => clk, Q => n74, 
                           QN => n_1883);
   MY_CLK_r_REG222_S4 : DFF_X1 port map( D => SIG_in(17), CK => clk, Q => n73, 
                           QN => n_1884);
   MY_CLK_r_REG221_S4 : DFF_X1 port map( D => SIG_in(16), CK => clk, Q => n72, 
                           QN => n_1885);
   MY_CLK_r_REG223_S4 : DFF_X1 port map( D => SIG_in(15), CK => clk, Q => n71, 
                           QN => n_1886);
   MY_CLK_r_REG204_S4 : DFF_X1 port map( D => SIG_in(14), CK => clk, Q => n70, 
                           QN => n_1887);
   MY_CLK_r_REG203_S4 : DFF_X1 port map( D => SIG_in(13), CK => clk, Q => n69, 
                           QN => n_1888);
   MY_CLK_r_REG225_S4 : DFF_X1 port map( D => SIG_in(12), CK => clk, Q => n68, 
                           QN => n_1889);
   MY_CLK_r_REG227_S4 : DFF_X1 port map( D => SIG_in(11), CK => clk, Q => n67, 
                           QN => n_1890);
   MY_CLK_r_REG243_S4 : DFF_X1 port map( D => SIG_in(10), CK => clk, Q => n66, 
                           QN => n_1891);
   MY_CLK_r_REG242_S4 : DFF_X1 port map( D => SIG_in(9), CK => clk, Q => n65, 
                           QN => n_1892);
   MY_CLK_r_REG241_S4 : DFF_X1 port map( D => SIG_in(8), CK => clk, Q => n64, 
                           QN => n_1893);
   MY_CLK_r_REG244_S4 : DFF_X1 port map( D => SIG_in(7), CK => clk, Q => n63, 
                           QN => n_1894);
   MY_CLK_r_REG245_S4 : DFF_X1 port map( D => SIG_in(6), CK => clk, Q => n62, 
                           QN => n_1895);
   MY_CLK_r_REG237_S4 : DFF_X1 port map( D => EXP_in(7), CK => clk, Q => n_1896
                           , QN => n86);
   MY_CLK_r_REG238_S4 : DFF_X1 port map( D => EXP_in(6), CK => clk, Q => n60, 
                           QN => n87);
   MY_CLK_r_REG236_S4 : DFF_X1 port map( D => EXP_in(5), CK => clk, Q => n59, 
                           QN => n85);
   MY_CLK_r_REG239_S4 : DFF_X1 port map( D => EXP_in(4), CK => clk, Q => n58, 
                           QN => n90);
   MY_CLK_r_REG235_S4 : DFF_X1 port map( D => EXP_in(3), CK => clk, Q => n57, 
                           QN => n_1897);
   MY_CLK_r_REG240_S4 : DFF_X1 port map( D => EXP_in(2), CK => clk, Q => n56, 
                           QN => n89);
   MY_CLK_r_REG247_S4 : DFF_X1 port map( D => EXP_in(1), CK => clk, Q => n55, 
                           QN => n_1898);
   MY_CLK_r_REG246_S4 : DFF_X1 port map( D => EXP_in(0), CK => clk, Q => n54, 
                           QN => n88);
   MY_CLK_r_REG211_S4 : DFF_X1 port map( D => SIG_in(27), CK => clk, Q => n53, 
                           QN => n_1899);
   MY_CLK_r_REG209_S4 : DFF_X1 port map( D => n25, CK => clk, Q => n51, QN => 
                           n97);
   U2 : NOR2_X1 port map( A1 => n11, A2 => n90, ZN => n94);
   U3 : AND2_X1 port map( A1 => n59, A2 => n58, ZN => n95);
   U4 : NAND3_X1 port map( A1 => n56, A2 => n57, A3 => n51, ZN => n11);
   U6 : XNOR2_X1 port map( A => n94, B => n85, ZN => EXP_out(5));
   U7 : NOR2_X1 port map( A1 => n16, A2 => n87, ZN => n93);
   U8 : XNOR2_X1 port map( A => n93, B => n86, ZN => EXP_out(7));
   U10 : NAND2_X1 port map( A1 => n98, A2 => n95, ZN => n16);
   U13 : AND3_X2 port map( A1 => n56, A2 => n57, A3 => n51, ZN => n98);
   U16 : AND3_X1 port map( A1 => EXP_in(1), A2 => SIG_in(27), A3 => EXP_in(0), 
                           ZN => n25);
   MY_CLK_r_REG210_S4 : DFF_X1 port map( D => SIG_in(27), CK => clk, Q => n52, 
                           QN => n_1900);

end SYN_FPnormalize;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPround_SIG_width28 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0));

end FPround_SIG_width28;

architecture SYN_FPround of FPround_SIG_width28 is

   component FPround_SIG_width28_DW01_inc_1
      port( A : in std_logic_vector (24 downto 0);  SUM : out std_logic_vector 
            (24 downto 0));
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, 
      N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, n30 : std_logic;

begin
   EXP_out <= ( EXP_in(7), EXP_in(6), EXP_in(5), EXP_in(4), EXP_in(3), 
      EXP_in(2), EXP_in(1), EXP_in(0) );
   
   U8 : MUX2_X1 port map( A => SIG_in(3), B => N2, S => SIG_in(2), Z => 
                           SIG_out(3));
   U9 : MUX2_X1 port map( A => SIG_in(4), B => N3, S => SIG_in(2), Z => 
                           SIG_out(4));
   U10 : MUX2_X1 port map( A => SIG_in(5), B => N4, S => SIG_in(2), Z => 
                           SIG_out(5));
   U11 : MUX2_X1 port map( A => SIG_in(6), B => N5, S => SIG_in(2), Z => 
                           SIG_out(6));
   U12 : MUX2_X1 port map( A => SIG_in(7), B => N6, S => SIG_in(2), Z => 
                           SIG_out(7));
   U13 : MUX2_X1 port map( A => SIG_in(8), B => N7, S => SIG_in(2), Z => 
                           SIG_out(8));
   U14 : MUX2_X1 port map( A => SIG_in(9), B => N8, S => SIG_in(2), Z => 
                           SIG_out(9));
   U15 : MUX2_X1 port map( A => SIG_in(10), B => N9, S => SIG_in(2), Z => 
                           SIG_out(10));
   U16 : MUX2_X1 port map( A => SIG_in(11), B => N10, S => SIG_in(2), Z => 
                           SIG_out(11));
   U17 : MUX2_X1 port map( A => SIG_in(12), B => N11, S => SIG_in(2), Z => 
                           SIG_out(12));
   U18 : MUX2_X1 port map( A => SIG_in(13), B => N12, S => SIG_in(2), Z => 
                           SIG_out(13));
   U19 : MUX2_X1 port map( A => SIG_in(14), B => N13, S => SIG_in(2), Z => 
                           SIG_out(14));
   U20 : MUX2_X1 port map( A => SIG_in(15), B => N14, S => SIG_in(2), Z => 
                           SIG_out(15));
   U21 : MUX2_X1 port map( A => SIG_in(16), B => N15, S => SIG_in(2), Z => 
                           SIG_out(16));
   U22 : MUX2_X1 port map( A => SIG_in(17), B => N16, S => SIG_in(2), Z => 
                           SIG_out(17));
   U23 : MUX2_X1 port map( A => SIG_in(18), B => N17, S => SIG_in(2), Z => 
                           SIG_out(18));
   U24 : MUX2_X1 port map( A => SIG_in(19), B => N18, S => SIG_in(2), Z => 
                           SIG_out(19));
   U25 : MUX2_X1 port map( A => SIG_in(20), B => N19, S => SIG_in(2), Z => 
                           SIG_out(20));
   U26 : MUX2_X1 port map( A => SIG_in(21), B => N20, S => SIG_in(2), Z => 
                           SIG_out(21));
   U27 : MUX2_X1 port map( A => SIG_in(22), B => N21, S => SIG_in(2), Z => 
                           SIG_out(22));
   U28 : MUX2_X1 port map( A => SIG_in(23), B => N22, S => SIG_in(2), Z => 
                           SIG_out(23));
   U29 : MUX2_X1 port map( A => SIG_in(24), B => N23, S => SIG_in(2), Z => 
                           SIG_out(24));
   U30 : MUX2_X1 port map( A => SIG_in(25), B => N24, S => SIG_in(2), Z => 
                           SIG_out(25));
   U31 : MUX2_X1 port map( A => SIG_in(26), B => N25, S => SIG_in(2), Z => 
                           SIG_out(26));
   n30 <= '0';
   U3 : AND2_X2 port map( A1 => N26, A2 => SIG_in(2), ZN => SIG_out(27));
   add_45 : FPround_SIG_width28_DW01_inc_1 port map( A(24) => n30, A(23) => 
                           SIG_in(26), A(22) => SIG_in(25), A(21) => SIG_in(24)
                           , A(20) => SIG_in(23), A(19) => SIG_in(22), A(18) =>
                           SIG_in(21), A(17) => SIG_in(20), A(16) => SIG_in(19)
                           , A(15) => SIG_in(18), A(14) => SIG_in(17), A(13) =>
                           SIG_in(16), A(12) => SIG_in(15), A(11) => SIG_in(14)
                           , A(10) => SIG_in(13), A(9) => SIG_in(12), A(8) => 
                           SIG_in(11), A(7) => SIG_in(10), A(6) => SIG_in(9), 
                           A(5) => SIG_in(8), A(4) => SIG_in(7), A(3) => 
                           SIG_in(6), A(2) => SIG_in(5), A(1) => SIG_in(4), 
                           A(0) => SIG_in(3), SUM(24) => N26, SUM(23) => N25, 
                           SUM(22) => N24, SUM(21) => N23, SUM(20) => N22, 
                           SUM(19) => N21, SUM(18) => N20, SUM(17) => N19, 
                           SUM(16) => N18, SUM(15) => N17, SUM(14) => N16, 
                           SUM(13) => N15, SUM(12) => N14, SUM(11) => N13, 
                           SUM(10) => N12, SUM(9) => N11, SUM(8) => N10, SUM(7)
                           => N9, SUM(6) => N8, SUM(5) => N7, SUM(4) => N6, 
                           SUM(3) => N5, SUM(2) => N4, SUM(1) => N3, SUM(0) => 
                           N2);

end SYN_FPround;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPnormalize_SIG_width28_0 is

   port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
         std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
         downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
         std_logic);

end FPnormalize_SIG_width28_0;

architecture SYN_FPnormalize of FPnormalize_SIG_width28_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n7, n8, n9, n11, n12, n14, n15, n17, n82, n83, n84, n133, 
      n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, 
      n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
      n170, n171, n172, n173, n174, n175, n176, n177, n178, n239, n240, n241, 
      n242, n243, n_1912, n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, 
      n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, 
      n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, 
      n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, 
      n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952 : std_logic;

begin
   
   U3 : XNOR2_X1 port map( A => n151, B => n14, ZN => EXP_out(6));
   U5 : XOR2_X1 port map( A => n133, B => n83, Z => EXP_out(0));
   U7 : NOR2_X1 port map( A1 => n243, A2 => n239, ZN => n4);
   U8 : XOR2_X1 port map( A => n136, B => n4, Z => EXP_out(1));
   U9 : NAND3_X1 port map( A1 => n136, A2 => n84, A3 => n133, ZN => n5);
   U10 : INV_X1 port map( A => n5, ZN => n8);
   U11 : XOR2_X1 port map( A => n139, B => n8, Z => EXP_out(2));
   U13 : NOR2_X1 port map( A1 => n241, A2 => n5, ZN => n7);
   U14 : XOR2_X1 port map( A => n142, B => n7, Z => EXP_out(3));
   U15 : NAND3_X1 port map( A1 => n142, A2 => n139, A3 => n8, ZN => n9);
   U16 : INV_X1 port map( A => n9, ZN => n12);
   U17 : XOR2_X1 port map( A => n145, B => n12, Z => EXP_out(4));
   U19 : NOR2_X1 port map( A1 => n242, A2 => n9, ZN => n11);
   U20 : XOR2_X1 port map( A => n148, B => n11, Z => EXP_out(5));
   U21 : NAND3_X1 port map( A1 => n148, A2 => n145, A3 => n12, ZN => n14);
   U23 : NOR2_X1 port map( A1 => n14, A2 => n240, ZN => n15);
   U24 : XOR2_X1 port map( A => n153, B => n15, Z => EXP_out(7));
   U29 : MUX2_X1 port map( A => n156, B => n157, S => n82, Z => SIG_out(3));
   U31 : MUX2_X1 port map( A => n158, B => n159, S => n83, Z => SIG_out(5));
   U32 : MUX2_X1 port map( A => n159, B => n160, S => n82, Z => SIG_out(6));
   U33 : MUX2_X1 port map( A => n160, B => n161, S => n83, Z => SIG_out(7));
   U34 : MUX2_X1 port map( A => n161, B => n162, S => n82, Z => SIG_out(8));
   U36 : MUX2_X1 port map( A => n163, B => n164, S => n83, Z => SIG_out(10));
   U37 : MUX2_X1 port map( A => n164, B => n165, S => n84, Z => SIG_out(11));
   U38 : MUX2_X1 port map( A => n165, B => n166, S => n84, Z => SIG_out(12));
   U39 : MUX2_X1 port map( A => n166, B => n167, S => n84, Z => SIG_out(13));
   U40 : MUX2_X1 port map( A => n167, B => n168, S => n84, Z => SIG_out(14));
   U41 : MUX2_X1 port map( A => n168, B => n169, S => n82, Z => SIG_out(15));
   U42 : MUX2_X1 port map( A => n169, B => n170, S => n84, Z => SIG_out(16));
   U43 : MUX2_X1 port map( A => n170, B => n171, S => n84, Z => SIG_out(17));
   U44 : MUX2_X1 port map( A => n171, B => n172, S => n82, Z => SIG_out(18));
   U45 : MUX2_X1 port map( A => n172, B => n173, S => n83, Z => SIG_out(19));
   U46 : MUX2_X1 port map( A => n173, B => n174, S => n82, Z => SIG_out(20));
   U47 : MUX2_X1 port map( A => n174, B => n175, S => n83, Z => SIG_out(21));
   U48 : MUX2_X1 port map( A => n175, B => n176, S => n82, Z => SIG_out(22));
   U49 : MUX2_X1 port map( A => n176, B => SIG_in(24), S => n83, Z => 
                           SIG_out(23));
   U50 : MUX2_X1 port map( A => SIG_in(24), B => n177, S => n82, Z => 
                           SIG_out(24));
   U51 : MUX2_X1 port map( A => n177, B => SIG_in(26), S => n82, Z => 
                           SIG_out(25));
   U52 : INV_X1 port map( A => SIG_in(26), ZN => n17);
   U53 : NAND2_X1 port map( A1 => n17, A2 => n243, ZN => SIG_out(26));
   U2 : BUF_X2 port map( A => n178, Z => n84);
   U6 : BUF_X1 port map( A => n178, Z => n83);
   U12 : BUF_X2 port map( A => n178, Z => n82);
   MY_CLK_r_REG234_S3 : DFF_X1 port map( D => SIG_in(27), CK => clk, Q => n178,
                           QN => n243);
   MY_CLK_r_REG233_S3 : DFF_X1 port map( D => SIG_in(25), CK => clk, Q => n177,
                           QN => n_1912);
   MY_CLK_r_REG229_S3 : DFF_X1 port map( D => SIG_in(23), CK => clk, Q => n176,
                           QN => n_1913);
   MY_CLK_r_REG231_S3 : DFF_X1 port map( D => SIG_in(22), CK => clk, Q => n175,
                           QN => n_1914);
   MY_CLK_r_REG230_S3 : DFF_X1 port map( D => SIG_in(21), CK => clk, Q => n174,
                           QN => n_1915);
   MY_CLK_r_REG232_S3 : DFF_X1 port map( D => SIG_in(20), CK => clk, Q => n173,
                           QN => n_1916);
   MY_CLK_r_REG249_S3 : DFF_X1 port map( D => SIG_in(19), CK => clk, Q => n172,
                           QN => n_1917);
   MY_CLK_r_REG252_S3 : DFF_X1 port map( D => SIG_in(18), CK => clk, Q => n171,
                           QN => n_1918);
   MY_CLK_r_REG251_S3 : DFF_X1 port map( D => SIG_in(17), CK => clk, Q => n170,
                           QN => n_1919);
   MY_CLK_r_REG250_S3 : DFF_X1 port map( D => SIG_in(16), CK => clk, Q => n169,
                           QN => n_1920);
   MY_CLK_r_REG228_S3 : DFF_X1 port map( D => SIG_in(15), CK => clk, Q => n168,
                           QN => n_1921);
   MY_CLK_r_REG202_S3 : DFF_X1 port map( D => SIG_in(14), CK => clk, Q => n167,
                           QN => n_1922);
   MY_CLK_r_REG224_S3 : DFF_X1 port map( D => SIG_in(13), CK => clk, Q => n166,
                           QN => n_1923);
   MY_CLK_r_REG226_S3 : DFF_X1 port map( D => SIG_in(12), CK => clk, Q => n165,
                           QN => n_1924);
   MY_CLK_r_REG255_S3 : DFF_X1 port map( D => SIG_in(11), CK => clk, Q => n164,
                           QN => n_1925);
   MY_CLK_r_REG254_S3 : DFF_X1 port map( D => SIG_in(10), CK => clk, Q => n163,
                           QN => n_1926);
   MY_CLK_r_REG253_S3 : DFF_X1 port map( D => SIG_in(9), CK => clk, Q => n162, 
                           QN => n_1927);
   MY_CLK_r_REG256_S3 : DFF_X1 port map( D => SIG_in(8), CK => clk, Q => n161, 
                           QN => n_1928);
   MY_CLK_r_REG258_S3 : DFF_X1 port map( D => SIG_in(7), CK => clk, Q => n160, 
                           QN => n_1929);
   MY_CLK_r_REG261_S3 : DFF_X1 port map( D => SIG_in(6), CK => clk, Q => n159, 
                           QN => n_1930);
   MY_CLK_r_REG264_S3 : DFF_X1 port map( D => SIG_in(5), CK => clk, Q => n158, 
                           QN => n_1931);
   MY_CLK_r_REG267_S3 : DFF_X1 port map( D => SIG_in(4), CK => clk, Q => n157, 
                           QN => n_1932);
   MY_CLK_r_REG271_S3 : DFF_X1 port map( D => SIG_in(3), CK => clk, Q => n156, 
                           QN => n_1933);
   MY_CLK_r_REG415_S3 : DFF_X1 port map( D => SIG_in(2), CK => clk, Q => n155, 
                           QN => n_1934);
   MY_CLK_r_REG386_S2 : DFF_X1 port map( D => EXP_in(7), CK => clk, Q => n154, 
                           QN => n_1935);
   MY_CLK_r_REG387_S3 : DFF_X1 port map( D => n154, CK => clk, Q => n153, QN =>
                           n_1936);
   MY_CLK_r_REG389_S2 : DFF_X1 port map( D => EXP_in(6), CK => clk, Q => n152, 
                           QN => n_1937);
   MY_CLK_r_REG390_S3 : DFF_X1 port map( D => n152, CK => clk, Q => n151, QN =>
                           n240);
   MY_CLK_r_REG392_S1 : DFF_X1 port map( D => EXP_in(5), CK => clk, Q => n150, 
                           QN => n_1938);
   MY_CLK_r_REG393_S2 : DFF_X1 port map( D => n150, CK => clk, Q => n149, QN =>
                           n_1939);
   MY_CLK_r_REG394_S3 : DFF_X1 port map( D => n149, CK => clk, Q => n148, QN =>
                           n_1940);
   MY_CLK_r_REG395_S1 : DFF_X1 port map( D => EXP_in(4), CK => clk, Q => n147, 
                           QN => n_1941);
   MY_CLK_r_REG396_S2 : DFF_X1 port map( D => n147, CK => clk, Q => n146, QN =>
                           n_1942);
   MY_CLK_r_REG397_S3 : DFF_X1 port map( D => n146, CK => clk, Q => n145, QN =>
                           n242);
   MY_CLK_r_REG398_S1 : DFF_X1 port map( D => EXP_in(3), CK => clk, Q => n144, 
                           QN => n_1943);
   MY_CLK_r_REG399_S2 : DFF_X1 port map( D => n144, CK => clk, Q => n143, QN =>
                           n_1944);
   MY_CLK_r_REG400_S3 : DFF_X1 port map( D => n143, CK => clk, Q => n142, QN =>
                           n_1945);
   MY_CLK_r_REG401_S1 : DFF_X1 port map( D => EXP_in(2), CK => clk, Q => n141, 
                           QN => n_1946);
   MY_CLK_r_REG402_S2 : DFF_X1 port map( D => n141, CK => clk, Q => n140, QN =>
                           n_1947);
   MY_CLK_r_REG403_S3 : DFF_X1 port map( D => n140, CK => clk, Q => n139, QN =>
                           n241);
   MY_CLK_r_REG404_S1 : DFF_X1 port map( D => EXP_in(1), CK => clk, Q => n138, 
                           QN => n_1948);
   MY_CLK_r_REG405_S2 : DFF_X1 port map( D => n138, CK => clk, Q => n137, QN =>
                           n_1949);
   MY_CLK_r_REG406_S3 : DFF_X1 port map( D => n137, CK => clk, Q => n136, QN =>
                           n_1950);
   MY_CLK_r_REG407_S1 : DFF_X1 port map( D => EXP_in(0), CK => clk, Q => n135, 
                           QN => n_1951);
   MY_CLK_r_REG408_S2 : DFF_X1 port map( D => n135, CK => clk, Q => n134, QN =>
                           n_1952);
   MY_CLK_r_REG409_S3 : DFF_X1 port map( D => n134, CK => clk, Q => n133, QN =>
                           n239);
   U4 : MUX2_X2 port map( A => n155, B => n156, S => n82, Z => SIG_out(2));
   U18 : MUX2_X1 port map( A => n158, B => n157, S => n243, Z => SIG_out(4));
   U22 : MUX2_X1 port map( A => n163, B => n162, S => n243, Z => SIG_out(9));

end SYN_FPnormalize;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity MBE is

   port( A, B : in std_logic_vector (31 downto 0);  C : out std_logic_vector 
         (63 downto 0);  clk : in std_logic);

end MBE;

architecture SYN_beh of MBE is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (63 downto 0);  Cout : out std_logic;  clk : 
            in std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_186
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR, clk : in 
            std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component HA_1
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_2
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_204
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);
   end component;
   
   component FA_205
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci : in std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component HA_4
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_5
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR, clk : in 
            std_logic);
   end component;
   
   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_288
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci, clk : in 
            std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_292
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component HA_7
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_8
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_306
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR, clk : in 
            std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_10
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_11
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_365
      port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_378
      port( A, B : in std_logic;  S, Co : out std_logic;  clk, Ci : in 
            std_logic);
   end component;
   
   component FA_379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_13
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_14
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_388
      port( A, Ci : in std_logic;  Co : out std_logic;  B_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_389
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR, clk : in 
            std_logic);
   end component;
   
   component FA_390
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR, clk : in 
            std_logic);
   end component;
   
   component FA_391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_16
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_17
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_19
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_20
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_477
      port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_479
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic
            );
   end component;
   
   component FA_480
      port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_482
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic
            );
   end component;
   
   component FA_483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_22
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_23
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_24
      port( B : in std_logic;  C, S_BAR : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_485
      port( B, Ci : in std_logic;  Co : out std_logic;  A_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_486
      port( A, Ci : in std_logic;  Co : out std_logic;  B_BAR : in std_logic;  
            S_BAR : out std_logic);
   end component;
   
   component FA_487
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_488
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_489
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_490
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_491
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_492
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_493
      port( A, B : in std_logic;  S, Co : out std_logic;  Ci_BAR : in std_logic
            );
   end component;
   
   component FA_494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_25
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_26
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_512
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_513
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_514
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_515
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_516
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_517
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_518
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_519
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_520
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_521
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_522
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_523
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_524
      port( A, B : in std_logic;  S, Co : out std_logic;  clk, Ci_BAR : in 
            std_logic);
   end component;
   
   component FA_525
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_526
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_527
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_528
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_529
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_530
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_531
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_532
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_533
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_534
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_535
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_536
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_28
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_29
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_539
      port( B, Ci : in std_logic;  S, Co : out std_logic;  A : in std_logic);
   end component;
   
   component FA_540
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_541
      port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_542
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_543
      port( A, Ci : in std_logic;  S, Co : out std_logic;  B_BAR : in std_logic
            );
   end component;
   
   component FA_544
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_545
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_546
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_547
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_548
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_549
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_550
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_551
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_552
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_553
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_554
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_555
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_556
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_557
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_558
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_559
      port( A, B, Ci : in std_logic;  S, Co : out std_logic;  clk : in 
            std_logic);
   end component;
   
   component FA_560
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_561
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_562
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_563
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_564
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_565
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_566
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_567
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_568
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_31
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_32
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_33
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_569
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_570
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_571
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_572
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_34
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_35
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_36
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_573
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_574
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_575
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_576
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_577
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_578
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_579
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_580
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_37
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_38
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_39
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_581
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_582
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_583
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_584
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_585
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_586
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_587
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_588
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_589
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_590
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_591
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_592
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_40
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_41
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_42
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component FA_593
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_594
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_595
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_596
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_597
      port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_598
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_599
      port( Ci : in std_logic;  S, Co : out std_logic;  B_BAR, A_BAR : in 
            std_logic);
   end component;
   
   component FA_600
      port( B, Ci : in std_logic;  S, Co : out std_logic;  A_BAR : in std_logic
            );
   end component;
   
   component FA_601
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_602
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_603
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_604
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_605
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_606
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_607
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component HA_43
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component HA_0
      port( A, B : in std_logic;  S, C : out std_logic);
   end component;
   
   component ENC_5
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  clk : in std_logic;  p_32_port, p_31_port, p_30_port, 
            p_29_port, p_28_port, p_27_port, p_26_port, p_25_port, p_24_port, 
            p_23_port, p_18_BAR, p_12_port, p_11_port, p_10_port, p_9_port, 
            p_8_port, p_6_port, p_3_port, p_1_port, p_0_port, p_17_BAR, 
            p_20_BAR, p_19_BAR, p_22_BAR, p_21_BAR, p_7_BAR, p_5_BAR, p_4_BAR, 
            p_2_BAR, p_14_BAR, p_13_BAR, p_16_BAR, p_15_BAR : out std_logic);
   end component;
   
   component ENC_6
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_7
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_8
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_9
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_10
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_11
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_12
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_13
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_14
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_15
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_16
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component ENC_0
      port( b : in std_logic_vector (2 downto 0);  A : in std_logic_vector (31 
            downto 0);  p : out std_logic_vector (32 downto 0);  clk : in 
            std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, n219, n220, q_0_0_32_port, 
      q_0_0_31_port, q_0_0_30_port, q_0_0_29_port, q_0_0_28_port, q_0_0_27_port
      , q_0_0_26_port, q_0_0_25_port, q_0_0_24_port, q_0_0_23_port, 
      q_0_0_22_port, q_0_0_21_port, q_0_0_20_port, q_0_0_19_port, q_0_0_18_port
      , q_0_0_17_port, q_0_0_16_port, q_0_0_15_port, q_0_0_14_port, 
      q_0_0_13_port, q_0_0_12_port, q_0_0_11_port, q_0_0_10_port, q_0_0_9_port,
      q_0_0_8_port, q_0_0_7_port, q_0_0_6_port, q_0_0_5_port, q_0_0_4_port, 
      q_0_0_3_port, q_0_0_2_port, q_0_0_1_port, q_0_0_0_port, q_0_8_42_port, 
      q_0_8_41_port, q_0_8_40_port, q_0_8_39_port, q_0_8_38_port, q_0_8_37_port
      , q_0_8_36_port, q_0_8_35_port, q_0_8_34_port, q_0_8_33_port, 
      q_0_8_32_port, q_0_8_31_port, q_0_8_30_port, q_0_8_29_port, q_0_8_28_port
      , q_0_8_27_port, q_0_8_26_port, q_0_8_25_port, q_0_8_24_port, 
      q_0_8_23_port, q_0_8_22_port, q_0_8_21_port, q_0_8_20_port, q_0_8_19_port
      , q_0_8_18_port, q_0_8_17_port, q_0_8_16_port, q_0_7_44_port, 
      q_0_7_43_port, q_0_7_42_port, q_0_7_41_port, q_0_7_40_port, q_0_7_39_port
      , q_0_7_38_port, q_0_7_37_port, q_0_7_36_port, q_0_7_35_port, 
      q_0_7_34_port, q_0_7_33_port, q_0_7_32_port, q_0_7_31_port, q_0_7_30_port
      , q_0_7_29_port, q_0_7_28_port, q_0_7_27_port, q_0_7_26_port, 
      q_0_7_25_port, q_0_7_24_port, q_0_7_23_port, q_0_7_22_port, q_0_7_21_port
      , q_0_7_20_port, q_0_7_19_port, q_0_7_18_port, q_0_7_17_port, 
      q_0_7_16_port, q_0_7_15_port, q_0_7_14_port, q_0_6_46_port, q_0_6_45_port
      , q_0_6_44_port, q_0_6_43_port, q_0_6_42_port, q_0_6_41_port, 
      q_0_6_40_port, q_0_6_39_port, q_0_6_38_port, q_0_6_37_port, q_0_6_36_port
      , q_0_6_35_port, q_0_6_34_port, q_0_6_33_port, q_0_6_32_port, 
      q_0_6_31_port, q_0_6_30_port, q_0_6_29_port, q_0_6_28_port, q_0_6_27_port
      , q_0_6_26_port, q_0_6_25_port, q_0_6_24_port, q_0_6_23_port, 
      q_0_6_22_port, q_0_6_21_port, q_0_6_20_port, q_0_6_19_port, q_0_6_18_port
      , q_0_6_17_port, q_0_6_16_port, q_0_6_15_port, q_0_6_14_port, 
      q_0_6_13_port, q_0_6_12_port, q_0_5_47_port, q_0_5_46_port, q_0_5_45_port
      , q_0_5_44_port, q_0_5_43_port, q_0_5_42_port, q_0_5_41_port, 
      q_0_5_40_port, q_0_5_39_port, q_0_5_38_port, q_0_5_37_port, q_0_5_36_port
      , q_0_5_35_port, q_0_5_34_port, q_0_5_33_port, q_0_5_32_port, 
      q_0_5_31_port, q_0_5_30_port, q_0_5_29_port, q_0_5_28_port, q_0_5_27_port
      , q_0_5_26_port, q_0_5_25_port, q_0_5_24_port, q_0_5_23_port, 
      q_0_5_22_port, q_0_5_21_port, q_0_5_20_port, q_0_5_19_port, q_0_5_18_port
      , q_0_5_17_port, q_0_5_16_port, q_0_5_15_port, q_0_5_14_port, 
      q_0_5_13_port, q_0_5_12_port, q_0_5_11_port, q_0_5_10_port, q_0_4_47_port
      , q_0_4_46_port, q_0_4_45_port, q_0_4_44_port, q_0_4_43_port, 
      q_0_4_42_port, q_0_4_41_port, q_0_4_40_port, q_0_4_39_port, q_0_4_38_port
      , q_0_4_37_port, q_0_4_36_port, q_0_4_35_port, q_0_4_34_port, 
      q_0_4_33_port, q_0_4_32_port, q_0_4_31_port, q_0_4_30_port, q_0_4_29_port
      , q_0_4_28_port, q_0_4_27_port, q_0_4_26_port, q_0_4_25_port, 
      q_0_4_24_port, q_0_4_23_port, q_0_4_22_port, q_0_4_21_port, q_0_4_20_port
      , q_0_4_19_port, q_0_4_18_port, q_0_4_17_port, q_0_4_16_port, 
      q_0_4_15_port, q_0_4_14_port, q_0_4_13_port, q_0_4_12_port, q_0_4_11_port
      , q_0_4_10_port, q_0_4_9_port, q_0_4_8_port, q_0_3_47_port, q_0_3_46_port
      , q_0_3_45_port, q_0_3_44_port, q_0_3_43_port, q_0_3_42_port, 
      q_0_3_41_port, q_0_3_40_port, q_0_3_39_port, q_0_3_38_port, q_0_3_37_port
      , q_0_3_36_port, q_0_3_35_port, q_0_3_34_port, q_0_3_33_port, 
      q_0_3_32_port, q_0_3_31_port, q_0_3_30_port, q_0_3_29_port, q_0_3_28_port
      , q_0_3_27_port, q_0_3_26_port, q_0_3_25_port, q_0_3_24_port, 
      q_0_3_23_port, q_0_3_22_port, q_0_3_21_port, q_0_3_20_port, q_0_3_19_port
      , q_0_3_18_port, q_0_3_17_port, q_0_3_16_port, q_0_3_15_port, 
      q_0_3_14_port, q_0_3_13_port, q_0_3_12_port, q_0_3_11_port, q_0_3_10_port
      , q_0_3_9_port, q_0_3_8_port, q_0_3_7_port, q_0_3_6_port, q_0_2_47_port, 
      q_0_2_46_port, q_0_2_45_port, q_0_2_44_port, q_0_2_43_port, q_0_2_42_port
      , q_0_2_41_port, q_0_2_40_port, q_0_2_39_port, q_0_2_38_port, 
      q_0_2_37_port, q_0_2_36_port, q_0_2_35_port, q_0_2_34_port, q_0_2_33_port
      , q_0_2_32_port, q_0_2_31_port, q_0_2_30_port, q_0_2_29_port, 
      q_0_2_28_port, q_0_2_27_port, q_0_2_26_port, q_0_2_25_port, q_0_2_24_port
      , q_0_2_23_port, q_0_2_22_port, q_0_2_21_port, q_0_2_20_port, 
      q_0_2_19_port, q_0_2_18_port, q_0_2_17_port, q_0_2_16_port, q_0_2_15_port
      , q_0_2_14_port, q_0_2_13_port, q_0_2_12_port, q_0_2_11_port, 
      q_0_2_10_port, q_0_2_9_port, q_0_2_8_port, q_0_2_7_port, q_0_2_6_port, 
      q_0_2_5_port, q_0_2_4_port, q_0_1_47_port, q_0_1_46_port, q_0_1_45_port, 
      q_0_1_44_port, q_0_1_43_port, q_0_1_42_port, q_0_1_41_port, q_0_1_40_port
      , q_0_1_39_port, q_0_1_38_port, q_0_1_37_port, q_0_1_36_port, 
      q_0_1_34_port, q_0_1_33_port, q_0_1_32_port, q_0_1_31_port, q_0_1_30_port
      , q_0_1_29_port, q_0_1_28_port, q_0_1_27_port, q_0_1_26_port, 
      q_0_1_25_port, q_0_1_24_port, q_0_1_23_port, q_0_1_21_port, q_0_1_20_port
      , q_0_1_19_port, q_0_1_18_port, q_0_1_17_port, q_0_1_16_port, 
      q_0_1_15_port, q_0_1_14_port, q_0_1_13_port, q_0_1_12_port, q_0_1_11_port
      , q_0_1_10_port, q_0_1_9_port, q_0_1_8_port, q_0_1_7_port, q_0_1_6_port, 
      q_0_1_5_port, q_0_1_4_port, q_0_1_3_port, q_0_1_2_port, q_0_12_35_port, 
      q_0_12_34_port, q_0_12_33_port, q_0_12_32_port, q_0_12_31_port, 
      q_0_12_30_port, q_0_12_29_port, q_0_12_28_port, q_0_12_27_port, 
      q_0_12_26_port, q_0_12_25_port, q_0_12_24_port, q_0_11_36_port, 
      q_0_11_35_port, q_0_11_34_port, q_0_11_33_port, q_0_11_32_port, 
      q_0_11_31_port, q_0_11_30_port, q_0_11_29_port, q_0_11_28_port, 
      q_0_11_27_port, q_0_11_26_port, q_0_11_25_port, q_0_11_24_port, 
      q_0_11_23_port, q_0_11_22_port, q_0_10_38_port, q_0_10_37_port, 
      q_0_10_36_port, q_0_10_35_port, q_0_10_34_port, q_0_10_33_port, 
      q_0_10_32_port, q_0_10_31_port, q_0_10_30_port, q_0_10_29_port, 
      q_0_10_28_port, q_0_10_27_port, q_0_10_26_port, q_0_10_25_port, 
      q_0_10_24_port, q_0_10_23_port, q_0_10_22_port, q_0_10_21_port, 
      q_0_10_20_port, q_0_9_40_port, q_0_9_39_port, q_0_9_38_port, 
      q_0_9_37_port, q_0_9_36_port, q_0_9_35_port, q_0_9_34_port, q_0_9_33_port
      , q_0_9_32_port, q_0_9_31_port, q_0_9_30_port, q_0_9_28_port, 
      q_0_9_27_port, q_0_9_26_port, q_0_9_25_port, q_0_9_24_port, q_0_9_23_port
      , q_0_9_22_port, q_0_9_21_port, q_0_9_20_port, q_0_9_19_port, 
      q_0_9_18_port, q_1_1_42_port, q_1_1_41_port, q_1_1_40_port, q_1_1_39_port
      , q_1_1_38_port, q_1_1_37_port, q_1_1_36_port, q_1_1_35_port, 
      q_1_1_34_port, q_1_1_33_port, q_1_1_32_port, q_1_1_31_port, q_1_1_30_port
      , q_1_1_29_port, q_1_1_28_port, q_1_1_26_port, q_1_1_25_port, 
      q_1_0_43_port, q_1_0_42_port, q_1_0_41_port, q_1_0_40_port, q_1_0_39_port
      , q_1_0_38_port, q_1_0_37_port, q_1_0_36_port, q_1_0_35_port, 
      q_1_0_34_port, q_1_0_33_port, q_1_0_32_port, q_1_0_31_port, q_1_0_30_port
      , q_1_0_27_port, q_1_0_26_port, q_1_0_25_port, q_1_0_24_port, 
      q_1_7_36_port, q_1_7_35_port, q_1_7_34_port, q_1_7_33_port, q_1_7_32_port
      , q_1_7_31_port, q_1_6_37_port, q_1_6_36_port, q_1_6_35_port, 
      q_1_6_34_port, q_1_6_33_port, q_1_6_32_port, q_1_6_31_port, q_1_6_30_port
      , q_1_5_38_port, q_1_5_37_port, q_1_5_36_port, q_1_5_35_port, 
      q_1_5_34_port, q_1_5_33_port, q_1_5_32_port, q_1_5_31_port, q_1_5_30_port
      , q_1_5_29_port, q_1_4_39_port, q_1_4_38_port, q_1_4_37_port, 
      q_1_4_36_port, q_1_4_35_port, q_1_4_34_port, q_1_4_33_port, q_1_4_32_port
      , q_1_4_31_port, q_1_4_30_port, q_1_4_29_port, q_1_4_28_port, 
      q_1_3_40_port, q_1_3_39_port, q_1_3_38_port, q_1_3_37_port, q_1_3_36_port
      , q_1_3_35_port, q_1_3_34_port, q_1_3_33_port, q_1_3_32_port, 
      q_1_3_31_port, q_1_3_30_port, q_1_3_28_port, q_1_3_27_port, q_1_2_41_port
      , q_1_2_40_port, q_1_2_39_port, q_1_2_38_port, q_1_2_37_port, 
      q_1_2_36_port, q_1_2_35_port, q_1_2_34_port, q_1_2_33_port, q_1_2_32_port
      , q_1_2_31_port, q_1_2_30_port, q_1_2_29_port, q_1_2_28_port, 
      q_1_2_26_port, q_2_2_47_port, q_2_2_46_port, q_2_2_45_port, q_2_2_44_port
      , q_2_2_43_port, q_2_2_42_port, q_2_2_41_port, q_2_2_40_port, 
      q_2_2_39_port, q_2_2_37_port, q_2_2_36_port, q_2_2_35_port, q_2_2_34_port
      , q_2_2_33_port, q_2_2_32_port, q_2_2_31_port, q_2_2_30_port, 
      q_2_2_29_port, q_2_2_28_port, q_2_2_27_port, q_2_2_26_port, q_2_2_25_port
      , q_2_2_24_port, q_2_2_23_port, q_2_2_22_port, q_2_2_21_port, 
      q_2_2_20_port, q_2_2_19_port, q_2_2_18_port, q_2_1_47_port, q_2_1_46_port
      , q_2_1_45_port, q_2_1_44_port, q_2_1_43_port, q_2_1_42_port, 
      q_2_1_41_port, q_2_1_40_port, q_2_1_39_port, q_2_1_38_port, q_2_1_37_port
      , q_2_1_36_port, q_2_1_35_port, q_2_1_34_port, q_2_1_33_port, 
      q_2_1_32_port, q_2_1_31_port, q_2_1_30_port, q_2_1_29_port, q_2_1_28_port
      , q_2_1_27_port, q_2_1_26_port, q_2_1_25_port, q_2_1_24_port, 
      q_2_1_23_port, q_2_1_22_port, q_2_1_21_port, q_2_1_20_port, q_2_1_19_port
      , q_2_1_18_port, q_2_1_17_port, q_2_0_47_port, q_2_0_46_port, 
      q_2_0_45_port, q_2_0_44_port, q_2_0_43_port, q_2_0_42_port, q_2_0_41_port
      , q_2_0_39_port, q_2_0_38_port, q_2_0_37_port, q_2_0_36_port, 
      q_2_0_35_port, q_2_0_33_port, q_2_0_32_port, q_2_0_31_port, q_2_0_30_port
      , q_2_0_29_port, q_2_0_28_port, q_2_0_27_port, q_2_0_26_port, 
      q_2_0_25_port, q_2_0_24_port, q_2_0_23_port, q_2_0_22_port, q_2_0_21_port
      , q_2_0_20_port, q_2_0_19_port, q_2_0_18_port, q_2_0_17_port, 
      q_2_0_16_port, q_2_7_30_port, q_2_7_28_port, q_2_7_27_port, q_2_7_26_port
      , q_2_7_25_port, q_2_7_24_port, q_2_7_23_port, q_2_6_31_port, 
      q_2_6_29_port, q_2_6_28_port, q_2_6_27_port, q_2_6_26_port, q_2_6_25_port
      , q_2_6_24_port, q_2_6_22_port, q_2_5_45_port, q_2_5_44_port, 
      q_2_5_43_port, q_2_5_42_port, q_2_5_41_port, q_2_5_40_port, q_2_5_39_port
      , q_2_5_38_port, q_2_5_37_port, q_2_5_36_port, q_2_5_35_port, 
      q_2_5_34_port, q_2_5_33_port, q_2_5_32_port, q_2_5_31_port, q_2_5_30_port
      , q_2_5_29_port, q_2_5_28_port, q_2_5_27_port, q_2_5_26_port, 
      q_2_5_25_port, q_2_5_24_port, q_2_5_23_port, q_2_5_22_port, q_2_5_21_port
      , q_2_4_46_port, q_2_4_45_port, q_2_4_44_port, q_2_4_43_port, 
      q_2_4_42_port, q_2_4_41_port, q_2_4_40_port, q_2_4_39_port, q_2_4_38_port
      , q_2_4_37_port, q_2_4_36_port, q_2_4_35_port, q_2_4_34_port, 
      q_2_4_33_port, q_2_4_32_port, q_2_4_31_port, q_2_4_30_port, q_2_4_29_port
      , q_2_4_28_port, q_2_4_27_port, q_2_4_26_port, q_2_4_25_port, 
      q_2_4_24_port, q_2_4_23_port, q_2_4_22_port, q_2_4_21_port, q_2_4_20_port
      , q_2_3_47_port, q_2_3_46_port, q_2_3_45_port, q_2_3_44_port, 
      q_2_3_43_port, q_2_3_42_port, q_2_3_41_port, q_2_3_40_port, q_2_3_39_port
      , q_2_3_38_port, q_2_3_37_port, q_2_3_36_port, q_2_3_35_port, 
      q_2_3_34_port, q_2_3_32_port, q_2_3_31_port, q_2_3_30_port, q_2_3_29_port
      , q_2_3_28_port, q_2_3_27_port, q_2_3_26_port, q_2_3_25_port, 
      q_2_3_24_port, q_2_3_23_port, q_2_3_22_port, q_2_3_21_port, q_2_3_20_port
      , q_2_3_19_port, q_3_3_47_port, q_3_3_46_port, q_3_3_45_port, 
      q_3_3_44_port, q_3_3_43_port, q_3_3_42_port, q_3_3_41_port, q_3_3_40_port
      , q_3_3_39_port, q_3_3_38_port, q_3_3_37_port, q_3_3_36_port, 
      q_3_3_35_port, q_3_3_34_port, q_3_3_33_port, q_3_3_32_port, q_3_3_31_port
      , q_3_3_30_port, q_3_3_28_port, q_3_3_27_port, q_3_3_26_port, 
      q_3_3_25_port, q_3_3_24_port, q_3_3_23_port, q_3_3_22_port, q_3_3_21_port
      , q_3_3_20_port, q_3_3_19_port, q_3_3_18_port, q_3_3_17_port, 
      q_3_3_16_port, q_3_3_15_port, q_3_3_14_port, q_3_3_13_port, q_3_2_47_port
      , q_3_2_46_port, q_3_2_45_port, q_3_2_44_port, q_3_2_42_port, 
      q_3_2_41_port, q_3_2_40_port, q_3_2_39_port, q_3_2_38_port, q_3_2_37_port
      , q_3_2_36_port, q_3_2_35_port, q_3_2_34_port, q_3_2_33_port, 
      q_3_2_32_port, q_3_2_29_port, q_3_2_28_port, q_3_2_27_port, q_3_2_26_port
      , q_3_2_25_port, q_3_2_24_port, q_3_2_23_port, q_3_2_22_port, 
      q_3_2_20_port, q_3_2_19_port, q_3_2_18_port, q_3_2_17_port, q_3_2_16_port
      , q_3_2_15_port, q_3_2_14_port, q_3_2_13_port, q_3_2_12_port, 
      q_3_1_47_port, q_3_1_46_port, q_3_1_45_port, q_3_1_43_port, q_3_1_42_port
      , q_3_1_41_port, q_3_1_40_port, q_3_1_39_port, q_3_1_38_port, 
      q_3_1_37_port, q_3_1_36_port, q_3_1_34_port, q_3_1_33_port, q_3_1_32_port
      , q_3_1_31_port, q_3_1_30_port, q_3_1_29_port, q_3_1_28_port, 
      q_3_1_27_port, q_3_1_26_port, q_3_1_25_port, q_3_1_24_port, q_3_1_23_port
      , q_3_1_22_port, q_3_1_21_port, q_3_1_20_port, q_3_1_19_port, 
      q_3_1_18_port, q_3_1_17_port, q_3_1_16_port, q_3_1_15_port, q_3_1_14_port
      , q_3_1_13_port, q_3_1_12_port, q_3_1_11_port, q_3_0_47_port, 
      q_3_0_46_port, q_3_0_45_port, q_3_0_44_port, q_3_0_42_port, q_3_0_41_port
      , q_3_0_40_port, q_3_0_39_port, q_3_0_38_port, q_3_0_37_port, 
      q_3_0_36_port, q_3_0_35_port, q_3_0_34_port, q_3_0_33_port, q_3_0_32_port
      , q_3_0_31_port, q_3_0_30_port, q_3_0_29_port, q_3_0_28_port, 
      q_3_0_27_port, q_3_0_26_port, q_3_0_25_port, q_3_0_24_port, q_3_0_22_port
      , q_3_0_21_port, q_3_0_20_port, q_3_0_19_port, q_3_0_18_port, 
      q_3_0_17_port, q_3_0_16_port, q_3_0_15_port, q_3_0_14_port, q_3_0_13_port
      , q_3_0_12_port, q_3_5_29_port, q_3_5_28_port, q_3_5_27_port, 
      q_3_5_26_port, q_3_5_25_port, q_3_5_24_port, q_3_5_23_port, q_3_5_22_port
      , q_3_5_21_port, q_3_5_20_port, q_3_5_19_port, q_3_5_18_port, 
      q_3_5_17_port, q_3_5_16_port, q_3_5_15_port, q_3_4_31_port, q_3_4_30_port
      , q_3_4_29_port, q_3_4_28_port, q_3_4_27_port, q_3_4_26_port, 
      q_3_4_25_port, q_3_4_24_port, q_3_4_23_port, q_3_4_22_port, q_3_4_21_port
      , q_3_4_20_port, q_3_4_19_port, q_3_4_18_port, q_3_4_17_port, 
      q_3_4_16_port, q_3_4_15_port, q_3_4_14_port, q_4_2_47_port, q_4_2_46_port
      , q_4_2_45_port, q_4_2_44_port, q_4_2_43_port, q_4_2_42_port, 
      q_4_2_41_port, q_4_2_40_port, q_4_2_39_port, q_4_2_38_port, q_4_2_37_port
      , q_4_2_36_port, q_4_2_35_port, q_4_2_34_port, q_4_2_33_port, 
      q_4_2_32_port, q_4_2_31_port, q_4_2_30_port, q_4_2_28_port, q_4_2_27_port
      , q_4_2_26_port, q_4_2_25_port, q_4_2_24_port, q_4_2_23_port, 
      q_4_2_22_port, q_4_2_21_port, q_4_2_20_port, q_4_2_19_port, q_4_2_18_port
      , q_4_2_17_port, q_4_2_16_port, q_4_2_15_port, q_4_2_14_port, 
      q_4_2_13_port, q_4_2_12_port, q_4_2_11_port, q_4_2_10_port, q_4_2_9_port,
      q_4_2_8_port, q_4_1_47_port, q_4_1_46_port, q_4_1_45_port, q_4_1_44_port,
      q_4_1_43_port, q_4_1_42_port, q_4_1_41_port, q_4_1_40_port, q_4_1_39_port
      , q_4_1_38_port, q_4_1_37_port, q_4_1_36_port, q_4_1_35_port, 
      q_4_1_34_port, q_4_1_33_port, q_4_1_32_port, q_4_1_31_port, q_4_1_30_port
      , q_4_1_29_port, q_4_1_28_port, q_4_1_26_port, q_4_1_25_port, 
      q_4_1_24_port, q_4_1_23_port, q_4_1_22_port, q_4_1_21_port, q_4_1_20_port
      , q_4_1_19_port, q_4_1_18_port, q_4_1_17_port, q_4_1_16_port, 
      q_4_1_15_port, q_4_1_14_port, q_4_1_13_port, q_4_1_12_port, q_4_1_11_port
      , q_4_1_10_port, q_4_1_9_port, q_4_1_8_port, q_4_1_7_port, q_4_0_47_port,
      q_4_0_46_port, q_4_0_45_port, q_4_0_44_port, q_4_0_43_port, q_4_0_42_port
      , q_4_0_41_port, q_4_0_40_port, q_4_0_39_port, q_4_0_38_port, 
      q_4_0_37_port, q_4_0_36_port, q_4_0_33_port, q_4_0_32_port, q_4_0_31_port
      , q_4_0_30_port, q_4_0_28_port, q_4_0_27_port, q_4_0_26_port, 
      q_4_0_25_port, q_4_0_24_port, q_4_0_23_port, q_4_0_22_port, q_4_0_21_port
      , q_4_0_20_port, q_4_0_19_port, q_4_0_18_port, q_4_0_17_port, 
      q_4_0_16_port, q_4_0_15_port, q_4_0_14_port, q_4_0_13_port, q_4_0_12_port
      , q_4_0_11_port, q_4_0_10_port, q_4_0_9_port, q_4_0_8_port, q_4_0_7_port,
      q_4_0_6_port, q_5_2_32_port, q_5_2_31_port, q_5_2_30_port, q_5_2_29_port,
      q_5_2_28_port, q_5_2_27_port, q_5_2_26_port, q_5_2_25_port, q_5_2_24_port
      , q_5_2_23_port, q_5_2_22_port, q_5_2_21_port, q_5_2_20_port, 
      q_5_2_19_port, q_5_2_18_port, q_5_2_17_port, q_5_2_16_port, q_5_2_15_port
      , q_5_2_14_port, q_5_2_13_port, q_5_2_12_port, q_5_2_11_port, 
      q_5_2_10_port, q_5_2_9_port, q_5_1_47_port, q_5_1_46_port, q_5_1_45_port,
      q_5_1_43_port, q_5_1_42_port, q_5_1_41_port, q_5_1_40_port, q_5_1_39_port
      , q_5_1_38_port, q_5_1_37_port, q_5_1_36_port, q_5_1_35_port, 
      q_5_1_34_port, q_5_1_33_port, q_5_1_32_port, q_5_1_31_port, q_5_1_30_port
      , q_5_1_29_port, q_5_1_27_port, q_5_1_26_port, q_5_1_25_port, 
      q_5_1_24_port, q_5_1_23_port, q_5_1_21_port, q_5_1_20_port, q_5_1_19_port
      , q_5_1_18_port, q_5_1_17_port, q_5_1_16_port, q_5_1_15_port, 
      q_5_1_14_port, q_5_1_13_port, q_5_1_12_port, q_5_1_11_port, q_5_1_10_port
      , q_5_1_9_port, q_5_1_8_port, q_5_1_6_port, q_5_1_5_port, q_5_0_47_port, 
      q_5_0_46_port, q_5_0_45_port, q_5_0_44_port, q_5_0_43_port, q_5_0_42_port
      , q_5_0_41_port, q_5_0_40_port, q_5_0_39_port, q_5_0_38_port, 
      q_5_0_37_port, q_5_0_36_port, q_5_0_35_port, q_5_0_34_port, q_5_0_33_port
      , q_5_0_32_port, q_5_0_31_port, q_5_0_30_port, q_5_0_29_port, 
      q_5_0_28_port, q_5_0_26_port, q_5_0_25_port, q_5_0_24_port, q_5_0_23_port
      , q_5_0_22_port, q_5_0_21_port, q_5_0_20_port, q_5_0_19_port, 
      q_5_0_18_port, q_5_0_17_port, q_5_0_16_port, q_5_0_15_port, q_5_0_14_port
      , q_5_0_13_port, q_5_0_12_port, q_5_0_11_port, q_5_0_10_port, 
      q_5_0_9_port, q_5_0_8_port, q_5_0_6_port, q_5_0_5_port, q_5_0_4_port, 
      q_6_1_47_port, q_6_1_46_port, q_6_1_45_port, q_6_1_44_port, q_6_1_43_port
      , q_6_1_42_port, q_6_1_41_port, q_6_1_40_port, q_6_1_39_port, 
      q_6_1_38_port, q_6_1_36_port, q_6_1_35_port, q_6_1_34_port, q_6_1_33_port
      , q_6_1_32_port, q_6_1_31_port, q_6_1_30_port, q_6_1_29_port, 
      q_6_1_28_port, q_6_1_27_port, q_6_1_26_port, q_6_1_25_port, q_6_1_24_port
      , q_6_1_23_port, q_6_1_22_port, q_6_1_21_port, q_6_1_20_port, 
      q_6_1_19_port, q_6_1_18_port, q_6_1_17_port, q_6_1_16_port, q_6_1_15_port
      , q_6_1_14_port, q_6_1_13_port, q_6_1_12_port, q_6_1_11_port, 
      q_6_1_10_port, q_6_1_9_port, q_6_1_8_port, q_6_1_7_port, q_6_1_6_port, 
      q_6_1_5_port, q_6_1_4_port, q_6_1_3_port, q_6_0_47_port, q_6_0_46_port, 
      q_6_0_45_port, q_6_0_44_port, q_6_0_43_port, q_6_0_42_port, q_6_0_41_port
      , q_6_0_40_port, q_6_0_39_port, q_6_0_38_port, q_6_0_37_port, 
      q_6_0_36_port, q_6_0_35_port, q_6_0_34_port, q_6_0_33_port, q_6_0_32_port
      , q_6_0_31_port, q_6_0_30_port, q_6_0_29_port, q_6_0_28_port, 
      q_6_0_27_port, q_6_0_26_port, q_6_0_25_port, q_6_0_24_port, q_6_0_23_port
      , q_6_0_22_port, q_6_0_21_port, q_6_0_20_port, q_6_0_19_port, 
      q_6_0_18_port, q_6_0_17_port, q_6_0_16_port, q_6_0_15_port, q_6_0_14_port
      , q_6_0_13_port, q_6_0_12_port, q_6_0_11_port, q_6_0_10_port, 
      q_6_0_9_port, q_6_0_8_port, q_6_0_7_port, q_6_0_6_port, q_6_0_5_port, 
      q_6_0_4_port, q_6_0_3_port, q_6_0_2_port, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n216, n218, net102736, net102737, net102738, net102739,
      net102740, net102741, net102742, net102743, net102744, net102745, 
      net102746, net102747, net102748, net102749, net102750, net102751, 
      net102752, net102753, net102754, net102755, net102756, net102757, 
      net102758, net102759, net102760, net102761, net102762, net102763, 
      net102764, net102765, net102766, net102767, net102768, net102769, 
      net102770, net102771, net102772, net102773, net102774, net102775, 
      net102776, net102777, net102778, net102779, net102780, net102781, 
      net102782, net102783, net102784, net102785, net102786, net102787, 
      net102788, net102789, net102790, net102791, net102792, net102793, 
      net102794, net102795, net102796, net102797, net102798, net102799, 
      net102800, net102801, net102802, net102803, net102804, net102805, 
      net102806, n227, n230, n233, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n373, 
      n374, n375, n376, n377, n379, n381, n382, n_2007, n_2008, n_2009, n_2010,
      n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, 
      n_2020, n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, 
      n_2029, n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, 
      n_2038, n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, 
      n_2047, n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, 
      n_2056, n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, 
      n_2065, n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, 
      n_2074, n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, 
      n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, 
      n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100 : 
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n182 <= '0';
   n183 <= '0';
   n184 <= '0';
   n185 <= '0';
   n186 <= '0';
   n187 <= '0';
   n188 <= '0';
   n189 <= '0';
   n190 <= '0';
   n191 <= '0';
   n192 <= '0';
   n193 <= '0';
   n194 <= '0';
   n195 <= '0';
   n196 <= '0';
   n197 <= '0';
   n198 <= '0';
   n199 <= '0';
   n200 <= '0';
   n201 <= '0';
   n202 <= '0';
   n203 <= '0';
   n204 <= '0';
   n205 <= '0';
   n206 <= '0';
   n207 <= '0';
   n208 <= '0';
   n209 <= '0';
   n210 <= '0';
   n211 <= '0';
   n212 <= '0';
   n213 <= '0';
   n220 <= '0';
   n219 <= '0';
   n218 <= '0';
   net102736 <= '0';
   net102737 <= '0';
   net102738 <= '0';
   net102739 <= '0';
   net102740 <= '0';
   net102741 <= '0';
   net102742 <= '0';
   net102743 <= '0';
   net102744 <= '0';
   net102745 <= '0';
   net102746 <= '0';
   net102747 <= '0';
   net102748 <= '0';
   net102749 <= '0';
   net102750 <= '0';
   net102751 <= '0';
   net102752 <= '0';
   net102753 <= '0';
   net102754 <= '0';
   net102755 <= '0';
   net102756 <= '0';
   net102757 <= '0';
   net102758 <= '0';
   net102759 <= '0';
   net102760 <= '0';
   net102761 <= '0';
   net102762 <= '0';
   net102763 <= '0';
   net102764 <= '0';
   net102765 <= '0';
   net102766 <= '0';
   net102767 <= '0';
   net102768 <= '0';
   net102769 <= '0';
   net102770 <= '0';
   net102771 <= '0';
   net102772 <= '0';
   net102773 <= '0';
   net102774 <= '0';
   net102775 <= '0';
   net102776 <= '0';
   net102777 <= '0';
   net102778 <= '0';
   net102779 <= '0';
   net102780 <= '0';
   net102781 <= '0';
   net102782 <= '0';
   net102783 <= '0';
   net102784 <= '0';
   net102785 <= '0';
   net102786 <= '0';
   net102787 <= '0';
   net102788 <= '0';
   net102789 <= '0';
   net102790 <= '0';
   net102791 <= '0';
   net102792 <= '0';
   net102793 <= '0';
   net102794 <= '0';
   net102795 <= '0';
   net102796 <= '0';
   net102797 <= '0';
   net102798 <= '0';
   net102799 <= '0';
   net102800 <= '0';
   net102801 <= '0';
   net102802 <= '0';
   net102803 <= '0';
   net102804 <= '0';
   net102805 <= '0';
   net102806 <= '0';
   U18 : INV_X1 port map( A => B(7), ZN => n227);
   U24 : INV_X1 port map( A => B(1), ZN => n233);
   U7 : BUF_X1 port map( A => A(23), Z => n382);
   U12 : INV_X1 port map( A => B(9), ZN => n216);
   U17 : BUF_X2 port map( A => B(23), Z => n379);
   U19 : INV_X1 port map( A => B(11), ZN => n230);
   encI_1 : ENC_0 port map( b(2) => B(1), b(1) => B(0), b(0) => X_Logic0_port, 
                           A(31) => n218, A(30) => n218, A(29) => n218, A(28) 
                           => n218, A(27) => n218, A(26) => n218, A(25) => n218
                           , A(24) => n218, A(23) => n381, A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), p(32) => 
                           q_0_0_32_port, p(31) => q_0_0_31_port, p(30) => 
                           q_0_0_30_port, p(29) => q_0_0_29_port, p(28) => 
                           q_0_0_28_port, p(27) => q_0_0_27_port, p(26) => 
                           q_0_0_26_port, p(25) => q_0_0_25_port, p(24) => 
                           q_0_0_24_port, p(23) => q_0_0_23_port, p(22) => 
                           q_0_0_22_port, p(21) => q_0_0_21_port, p(20) => 
                           q_0_0_20_port, p(19) => q_0_0_19_port, p(18) => 
                           q_0_0_18_port, p(17) => q_0_0_17_port, p(16) => 
                           q_0_0_16_port, p(15) => q_0_0_15_port, p(14) => 
                           q_0_0_14_port, p(13) => q_0_0_13_port, p(12) => 
                           q_0_0_12_port, p(11) => q_0_0_11_port, p(10) => 
                           q_0_0_10_port, p(9) => q_0_0_9_port, p(8) => 
                           q_0_0_8_port, p(7) => q_0_0_7_port, p(6) => 
                           q_0_0_6_port, p(5) => q_0_0_5_port, p(4) => 
                           q_0_0_4_port, p(3) => q_0_0_3_port, p(2) => 
                           q_0_0_2_port, p(1) => q_0_0_1_port, p(0) => 
                           q_0_0_0_port, clk => clk);
   encI_2 : ENC_16 port map( b(2) => B(3), b(1) => B(2), b(0) => B(1), A(31) =>
                           n218, A(30) => n218, A(29) => n218, A(28) => n218, 
                           A(27) => n218, A(26) => n218, A(25) => n218, A(24) 
                           => n218, A(23) => n382, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_34_port, p(31)
                           => q_0_1_33_port, p(30) => q_0_1_32_port, p(29) => 
                           q_0_1_31_port, p(28) => q_0_1_30_port, p(27) => 
                           q_0_1_29_port, p(26) => q_0_1_28_port, p(25) => 
                           q_0_1_27_port, p(24) => q_0_1_26_port, p(23) => 
                           q_0_1_25_port, p(22) => q_0_1_24_port, p(21) => 
                           q_0_1_23_port, p(20) => n362, p(19) => q_0_1_21_port
                           , p(18) => q_0_1_20_port, p(17) => q_0_1_19_port, 
                           p(16) => q_0_1_18_port, p(15) => q_0_1_17_port, 
                           p(14) => q_0_1_16_port, p(13) => q_0_1_15_port, 
                           p(12) => q_0_1_14_port, p(11) => q_0_1_13_port, 
                           p(10) => q_0_1_12_port, p(9) => q_0_1_11_port, p(8) 
                           => q_0_1_10_port, p(7) => q_0_1_9_port, p(6) => 
                           q_0_1_8_port, p(5) => q_0_1_7_port, p(4) => 
                           q_0_1_6_port, p(3) => q_0_1_5_port, p(2) => 
                           q_0_1_4_port, p(1) => q_0_1_3_port, p(0) => 
                           q_0_1_2_port, clk => clk);
   encI_3 : ENC_15 port map( b(2) => B(5), b(1) => B(4), b(0) => B(3), A(31) =>
                           n218, A(30) => n218, A(29) => n218, A(28) => n218, 
                           A(27) => n218, A(26) => n218, A(25) => n218, A(24) 
                           => n218, A(23) => n382, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_36_port, p(31)
                           => q_0_2_35_port, p(30) => q_0_2_34_port, p(29) => 
                           q_0_2_33_port, p(28) => q_0_2_32_port, p(27) => 
                           q_0_2_31_port, p(26) => q_0_2_30_port, p(25) => 
                           q_0_2_29_port, p(24) => q_0_2_28_port, p(23) => 
                           q_0_2_27_port, p(22) => q_0_2_26_port, p(21) => 
                           q_0_2_25_port, p(20) => q_0_2_24_port, p(19) => 
                           q_0_2_23_port, p(18) => q_0_2_22_port, p(17) => 
                           q_0_2_21_port, p(16) => q_0_2_20_port, p(15) => 
                           q_0_2_19_port, p(14) => q_0_2_18_port, p(13) => 
                           q_0_2_17_port, p(12) => q_0_2_16_port, p(11) => 
                           q_0_2_15_port, p(10) => q_0_2_14_port, p(9) => 
                           q_0_2_13_port, p(8) => q_0_2_12_port, p(7) => 
                           q_0_2_11_port, p(6) => q_0_2_10_port, p(5) => 
                           q_0_2_9_port, p(4) => q_0_2_8_port, p(3) => 
                           q_0_2_7_port, p(2) => q_0_2_6_port, p(1) => 
                           q_0_2_5_port, p(0) => q_0_2_4_port, clk => clk);
   encI_4 : ENC_14 port map( b(2) => B(7), b(1) => B(6), b(0) => B(5), A(31) =>
                           n218, A(30) => n218, A(29) => n218, A(28) => n218, 
                           A(27) => n218, A(26) => n218, A(25) => n218, A(24) 
                           => n218, A(23) => n381, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_38_port, p(31)
                           => q_0_1_37_port, p(30) => q_0_2_36_port, p(29) => 
                           q_0_3_35_port, p(28) => q_0_3_34_port, p(27) => 
                           q_0_3_33_port, p(26) => q_0_3_32_port, p(25) => 
                           q_0_3_31_port, p(24) => q_0_3_30_port, p(23) => 
                           q_0_3_29_port, p(22) => q_0_3_28_port, p(21) => 
                           q_0_3_27_port, p(20) => q_0_3_26_port, p(19) => 
                           q_0_3_25_port, p(18) => q_0_3_24_port, p(17) => 
                           q_0_3_23_port, p(16) => q_0_3_22_port, p(15) => 
                           q_0_3_21_port, p(14) => q_0_3_20_port, p(13) => 
                           q_0_3_19_port, p(12) => q_0_3_18_port, p(11) => 
                           q_0_3_17_port, p(10) => q_0_3_16_port, p(9) => 
                           q_0_3_15_port, p(8) => q_0_3_14_port, p(7) => 
                           q_0_3_13_port, p(6) => q_0_3_12_port, p(5) => 
                           q_0_3_11_port, p(4) => q_0_3_10_port, p(3) => 
                           q_0_3_9_port, p(2) => q_0_3_8_port, p(1) => 
                           q_0_3_7_port, p(0) => q_0_3_6_port, clk => clk);
   encI_5 : ENC_13 port map( b(2) => B(9), b(1) => B(8), b(0) => B(7), A(31) =>
                           n218, A(30) => n218, A(29) => n218, A(28) => n218, 
                           A(27) => n218, A(26) => n218, A(25) => n218, A(24) 
                           => n218, A(23) => n382, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_40_port, p(31)
                           => q_0_1_39_port, p(30) => q_0_2_38_port, p(29) => 
                           q_0_2_37_port, p(28) => q_0_3_36_port, p(27) => 
                           q_0_4_35_port, p(26) => q_0_4_34_port, p(25) => 
                           q_0_4_33_port, p(24) => q_0_4_32_port, p(23) => 
                           q_0_4_31_port, p(22) => q_0_4_30_port, p(21) => 
                           q_0_4_29_port, p(20) => q_0_4_28_port, p(19) => 
                           q_0_4_27_port, p(18) => q_0_4_26_port, p(17) => 
                           q_0_4_25_port, p(16) => q_0_4_24_port, p(15) => 
                           q_0_4_23_port, p(14) => q_0_4_22_port, p(13) => 
                           q_0_4_21_port, p(12) => q_0_4_20_port, p(11) => 
                           q_0_4_19_port, p(10) => q_0_4_18_port, p(9) => 
                           q_0_4_17_port, p(8) => q_0_4_16_port, p(7) => 
                           q_0_4_15_port, p(6) => q_0_4_14_port, p(5) => 
                           q_0_4_13_port, p(4) => q_0_4_12_port, p(3) => 
                           q_0_4_11_port, p(2) => q_0_4_10_port, p(1) => 
                           q_0_4_9_port, p(0) => q_0_4_8_port, clk => clk);
   encI_6 : ENC_12 port map( b(2) => B(11), b(1) => B(10), b(0) => B(9), A(31) 
                           => n218, A(30) => n218, A(29) => n218, A(28) => n218
                           , A(27) => n218, A(26) => n218, A(25) => n218, A(24)
                           => n218, A(23) => n381, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_42_port, p(31)
                           => q_0_1_41_port, p(30) => q_0_2_40_port, p(29) => 
                           q_0_2_39_port, p(28) => q_0_3_38_port, p(27) => 
                           q_0_3_37_port, p(26) => q_0_4_36_port, p(25) => 
                           q_0_5_35_port, p(24) => q_0_5_34_port, p(23) => 
                           q_0_5_33_port, p(22) => q_0_5_32_port, p(21) => 
                           q_0_5_31_port, p(20) => q_0_5_30_port, p(19) => 
                           q_0_5_29_port, p(18) => q_0_5_28_port, p(17) => 
                           q_0_5_27_port, p(16) => q_0_5_26_port, p(15) => 
                           q_0_5_25_port, p(14) => q_0_5_24_port, p(13) => 
                           q_0_5_23_port, p(12) => q_0_5_22_port, p(11) => 
                           q_0_5_21_port, p(10) => q_0_5_20_port, p(9) => 
                           q_0_5_19_port, p(8) => q_0_5_18_port, p(7) => 
                           q_0_5_17_port, p(6) => q_0_5_16_port, p(5) => 
                           q_0_5_15_port, p(4) => q_0_5_14_port, p(3) => 
                           q_0_5_13_port, p(2) => q_0_5_12_port, p(1) => 
                           q_0_5_11_port, p(0) => q_0_5_10_port, clk => clk);
   encI_7 : ENC_11 port map( b(2) => B(13), b(1) => B(12), b(0) => B(11), A(31)
                           => n218, A(30) => n218, A(29) => n218, A(28) => n218
                           , A(27) => n218, A(26) => n218, A(25) => n218, A(24)
                           => n218, A(23) => n381, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_44_port, p(31)
                           => q_0_1_43_port, p(30) => q_0_2_42_port, p(29) => 
                           q_0_2_41_port, p(28) => q_0_3_40_port, p(27) => 
                           q_0_3_39_port, p(26) => q_0_4_38_port, p(25) => 
                           q_0_4_37_port, p(24) => q_0_5_36_port, p(23) => 
                           q_0_6_35_port, p(22) => q_0_6_34_port, p(21) => 
                           q_0_6_33_port, p(20) => q_0_6_32_port, p(19) => 
                           q_0_6_31_port, p(18) => q_0_6_30_port, p(17) => 
                           q_0_6_29_port, p(16) => q_0_6_28_port, p(15) => 
                           q_0_6_27_port, p(14) => q_0_6_26_port, p(13) => 
                           q_0_6_25_port, p(12) => q_0_6_24_port, p(11) => 
                           q_0_6_23_port, p(10) => q_0_6_22_port, p(9) => 
                           q_0_6_21_port, p(8) => q_0_6_20_port, p(7) => 
                           q_0_6_19_port, p(6) => q_0_6_18_port, p(5) => 
                           q_0_6_17_port, p(4) => q_0_6_16_port, p(3) => 
                           q_0_6_15_port, p(2) => q_0_6_14_port, p(1) => 
                           q_0_6_13_port, p(0) => q_0_6_12_port, clk => clk);
   encI_8 : ENC_10 port map( b(2) => B(15), b(1) => B(14), b(0) => B(13), A(31)
                           => n218, A(30) => n218, A(29) => n218, A(28) => n218
                           , A(27) => n218, A(26) => n218, A(25) => n218, A(24)
                           => n218, A(23) => n381, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => q_0_1_46_port, p(31)
                           => q_0_1_45_port, p(30) => q_0_2_44_port, p(29) => 
                           q_0_2_43_port, p(28) => q_0_3_42_port, p(27) => 
                           q_0_3_41_port, p(26) => q_0_4_40_port, p(25) => 
                           q_0_4_39_port, p(24) => q_0_5_38_port, p(23) => 
                           q_0_5_37_port, p(22) => q_0_6_36_port, p(21) => 
                           q_0_7_35_port, p(20) => q_0_7_34_port, p(19) => 
                           q_0_7_33_port, p(18) => q_0_7_32_port, p(17) => 
                           q_0_7_31_port, p(16) => q_0_7_30_port, p(15) => 
                           q_0_7_29_port, p(14) => q_0_7_28_port, p(13) => 
                           q_0_7_27_port, p(12) => q_0_7_26_port, p(11) => 
                           q_0_7_25_port, p(10) => q_0_7_24_port, p(9) => 
                           q_0_7_23_port, p(8) => q_0_7_22_port, p(7) => 
                           q_0_7_21_port, p(6) => q_0_7_20_port, p(5) => 
                           q_0_7_19_port, p(4) => q_0_7_18_port, p(3) => 
                           q_0_7_17_port, p(2) => q_0_7_16_port, p(1) => 
                           q_0_7_15_port, p(0) => q_0_7_14_port, clk => clk);
   encI_9 : ENC_9 port map( b(2) => B(17), b(1) => B(16), b(0) => B(15), A(31) 
                           => n218, A(30) => n218, A(29) => n218, A(28) => n218
                           , A(27) => n218, A(26) => n218, A(25) => n218, A(24)
                           => n218, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2007, p(31) => 
                           q_0_1_47_port, p(30) => q_0_2_46_port, p(29) => 
                           q_0_2_45_port, p(28) => q_0_3_44_port, p(27) => 
                           q_0_3_43_port, p(26) => q_0_4_42_port, p(25) => 
                           q_0_4_41_port, p(24) => q_0_5_40_port, p(23) => 
                           q_0_5_39_port, p(22) => q_0_6_38_port, p(21) => 
                           q_0_6_37_port, p(20) => q_0_7_36_port, p(19) => 
                           q_0_8_35_port, p(18) => q_0_8_34_port, p(17) => 
                           q_0_8_33_port, p(16) => q_0_8_32_port, p(15) => 
                           q_0_8_31_port, p(14) => q_0_8_30_port, p(13) => 
                           q_0_8_29_port, p(12) => q_0_8_28_port, p(11) => 
                           q_0_8_27_port, p(10) => q_0_8_26_port, p(9) => 
                           q_0_8_25_port, p(8) => q_0_8_24_port, p(7) => 
                           q_0_8_23_port, p(6) => q_0_8_22_port, p(5) => 
                           q_0_8_21_port, p(4) => q_0_8_20_port, p(3) => 
                           q_0_8_19_port, p(2) => q_0_8_18_port, p(1) => 
                           q_0_8_17_port, p(0) => q_0_8_16_port, clk => clk);
   encI_10 : ENC_8 port map( b(2) => B(19), b(1) => B(18), b(0) => B(17), A(31)
                           => n218, A(30) => n218, A(29) => n218, A(28) => n218
                           , A(27) => n218, A(26) => n218, A(25) => n218, A(24)
                           => n218, A(23) => n381, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2008, p(31) => 
                           n_2009, p(30) => n_2010, p(29) => q_0_2_47_port, 
                           p(28) => q_0_3_46_port, p(27) => q_0_3_45_port, 
                           p(26) => q_0_4_44_port, p(25) => q_0_4_43_port, 
                           p(24) => q_0_5_42_port, p(23) => q_0_5_41_port, 
                           p(22) => q_0_6_40_port, p(21) => q_0_6_39_port, 
                           p(20) => q_0_7_38_port, p(19) => q_0_7_37_port, 
                           p(18) => q_0_8_36_port, p(17) => q_0_9_35_port, 
                           p(16) => q_0_9_34_port, p(15) => q_0_9_33_port, 
                           p(14) => q_0_9_32_port, p(13) => q_0_9_31_port, 
                           p(12) => q_0_9_30_port, p(11) => n361, p(10) => 
                           q_0_9_28_port, p(9) => q_0_9_27_port, p(8) => 
                           q_0_9_26_port, p(7) => q_0_9_25_port, p(6) => 
                           q_0_9_24_port, p(5) => q_0_9_23_port, p(4) => 
                           q_0_9_22_port, p(3) => q_0_9_21_port, p(2) => 
                           q_0_9_20_port, p(1) => q_0_9_19_port, p(0) => 
                           q_0_9_18_port, clk => clk);
   encI_11 : ENC_7 port map( b(2) => B(21), b(1) => B(20), b(0) => B(19), A(31)
                           => n218, A(30) => n218, A(29) => n218, A(28) => n218
                           , A(27) => n218, A(26) => n218, A(25) => n218, A(24)
                           => n218, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2011, p(31) => 
                           n_2012, p(30) => n_2013, p(29) => n_2014, p(28) => 
                           n_2015, p(27) => q_0_3_47_port, p(26) => 
                           q_0_4_46_port, p(25) => q_0_4_45_port, p(24) => 
                           q_0_5_44_port, p(23) => q_0_5_43_port, p(22) => 
                           q_0_6_42_port, p(21) => q_0_6_41_port, p(20) => 
                           q_0_7_40_port, p(19) => q_0_7_39_port, p(18) => 
                           q_0_8_38_port, p(17) => q_0_8_37_port, p(16) => 
                           q_0_9_36_port, p(15) => q_0_10_35_port, p(14) => 
                           q_0_10_34_port, p(13) => q_0_10_33_port, p(12) => 
                           q_0_10_32_port, p(11) => q_0_10_31_port, p(10) => 
                           q_0_10_30_port, p(9) => q_0_10_29_port, p(8) => 
                           q_0_10_28_port, p(7) => q_0_10_27_port, p(6) => 
                           q_0_10_26_port, p(5) => q_0_10_25_port, p(4) => 
                           q_0_10_24_port, p(3) => q_0_10_23_port, p(2) => 
                           q_0_10_22_port, p(1) => q_0_10_21_port, p(0) => 
                           q_0_10_20_port, clk => clk);
   encI_12 : ENC_6 port map( b(2) => B(23), b(1) => B(22), b(0) => B(21), A(31)
                           => n218, A(30) => n218, A(29) => n218, A(28) => n218
                           , A(27) => n218, A(26) => n218, A(25) => n218, A(24)
                           => n218, A(23) => n381, A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), p(32) => n_2016, p(31) => 
                           n_2017, p(30) => n_2018, p(29) => n_2019, p(28) => 
                           n_2020, p(27) => n_2021, p(26) => n_2022, p(25) => 
                           q_0_4_47_port, p(24) => q_0_5_46_port, p(23) => 
                           q_0_5_45_port, p(22) => q_0_6_44_port, p(21) => 
                           q_0_6_43_port, p(20) => q_0_7_42_port, p(19) => 
                           q_0_7_41_port, p(18) => q_0_8_40_port, p(17) => 
                           q_0_8_39_port, p(16) => q_0_9_38_port, p(15) => 
                           q_0_9_37_port, p(14) => q_0_10_36_port, p(13) => 
                           q_0_11_35_port, p(12) => q_0_11_34_port, p(11) => 
                           q_0_11_33_port, p(10) => q_0_11_32_port, p(9) => 
                           q_0_11_31_port, p(8) => q_0_11_30_port, p(7) => 
                           q_0_11_29_port, p(6) => q_0_11_28_port, p(5) => 
                           q_0_11_27_port, p(4) => q_0_11_26_port, p(3) => 
                           q_0_11_25_port, p(2) => q_0_11_24_port, p(1) => 
                           q_0_11_23_port, p(0) => q_0_11_22_port, clk => clk);
   encI_13 : ENC_5 port map( b(2) => n219, b(1) => n220, b(0) => n379, A(31) =>
                           n218, A(30) => n218, A(29) => n218, A(28) => n218, 
                           A(27) => n218, A(26) => n218, A(25) => n218, A(24) 
                           => n218, A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), clk => clk, p_32_port => 
                           n_2023, p_31_port => n_2024, p_30_port => n_2025, 
                           p_29_port => n_2026, p_28_port => n_2027, p_27_port 
                           => n_2028, p_26_port => n_2029, p_25_port => n_2030,
                           p_24_port => n_2031, p_23_port => q_0_5_47_port, 
                           p_18_BAR => q_0_8_42_port, p_12_port => 
                           q_0_11_36_port, p_11_port => q_0_12_35_port, 
                           p_10_port => q_0_12_34_port, p_9_port => 
                           q_0_12_33_port, p_8_port => q_0_12_32_port, p_6_port
                           => q_0_12_30_port, p_3_port => q_0_12_27_port, 
                           p_1_port => q_0_12_25_port, p_0_port => 
                           q_0_12_24_port, p_17_BAR => q_0_8_41_port, p_20_BAR 
                           => q_0_7_44_port, p_19_BAR => q_0_7_43_port, 
                           p_22_BAR => q_0_6_46_port, p_21_BAR => q_0_6_45_port
                           , p_7_BAR => q_0_12_31_port, p_5_BAR => 
                           q_0_12_29_port, p_4_BAR => q_0_12_28_port, p_2_BAR 
                           => q_0_12_26_port, p_14_BAR => q_0_10_38_port, 
                           p_13_BAR => q_0_10_37_port, p_16_BAR => 
                           q_0_9_40_port, p_15_BAR => q_0_9_39_port);
   HA_R_0_0_24 : HA_0 port map( A => q_0_0_24_port, B => q_0_1_24_port, S => 
                           q_1_0_24_port, C => q_1_1_25_port);
   HA_R_0_0_25 : HA_43 port map( A => q_0_0_25_port, B => q_0_1_25_port, S => 
                           q_1_0_25_port, C => q_1_1_26_port);
   FA_C_0_0_26 : FA_0 port map( A => q_0_0_26_port, B => q_0_1_26_port, Ci => 
                           q_0_2_26_port, S => q_1_0_26_port, Co => n351);
   FA_C_0_0_27 : FA_607 port map( A => q_0_0_27_port, B => q_0_1_27_port, Ci =>
                           q_0_2_27_port, S => q_1_0_27_port, Co => 
                           q_1_1_28_port);
   FA_C_0_0_28 : FA_606 port map( A => q_0_0_28_port, B => q_0_1_28_port, Ci =>
                           q_0_2_28_port, S => n348, Co => q_1_1_29_port);
   FA_C_0_0_29 : FA_605 port map( A => q_0_0_29_port, B => q_0_1_29_port, Ci =>
                           q_0_2_29_port, S => n352, Co => q_1_1_30_port);
   FA_C_0_0_30 : FA_604 port map( A => q_0_0_30_port, B => q_0_1_30_port, Ci =>
                           q_0_2_30_port, S => q_1_0_30_port, Co => 
                           q_1_1_31_port);
   FA_C_0_0_31 : FA_603 port map( A => q_0_0_31_port, B => q_0_1_31_port, Ci =>
                           q_0_2_31_port, S => q_1_0_31_port, Co => 
                           q_1_1_32_port);
   FA_C_0_0_32 : FA_602 port map( A => q_0_0_32_port, B => q_0_1_32_port, Ci =>
                           q_0_2_32_port, S => q_1_0_32_port, Co => 
                           q_1_1_33_port);
   FA_C_0_0_33 : FA_601 port map( A => B(1), B => q_0_1_33_port, Ci => 
                           q_0_2_33_port, S => q_1_0_33_port, Co => 
                           q_1_1_34_port);
   FA_C_0_0_34 : FA_600 port map( B => q_0_1_34_port, Ci => q_0_2_34_port, S =>
                           q_1_0_34_port, Co => q_1_1_35_port, A_BAR => n233);
   FA_C_0_0_35 : FA_599 port map( Ci => q_0_2_35_port, S => q_1_0_35_port, Co 
                           => q_1_1_36_port, B_BAR => B(3), A_BAR => B(1));
   FA_C_0_0_36 : FA_598 port map( A => X_Logic1_port, B => q_0_1_36_port, Ci =>
                           q_0_2_36_port, S => q_1_0_36_port, Co => 
                           q_1_1_37_port);
   FA_C_0_0_37 : FA_597 port map( B => q_0_1_37_port, Ci => q_0_2_37_port, S =>
                           q_1_0_37_port, Co => q_1_1_38_port, A_BAR => B(5));
   FA_C_0_0_38 : FA_596 port map( A => X_Logic1_port, B => q_0_1_38_port, Ci =>
                           q_0_2_38_port, S => q_1_0_38_port, Co => 
                           q_1_1_39_port);
   FA_C_0_0_39 : FA_595 port map( A => n227, B => q_0_1_39_port, Ci => 
                           q_0_2_39_port, S => q_1_0_39_port, Co => 
                           q_1_1_40_port);
   FA_C_0_0_40 : FA_594 port map( A => X_Logic1_port, B => q_0_1_40_port, Ci =>
                           q_0_2_40_port, S => q_1_0_40_port, Co => 
                           q_1_1_41_port);
   FA_C_0_0_41 : FA_593 port map( A => n216, B => q_0_1_41_port, Ci => 
                           q_0_2_41_port, S => q_1_0_41_port, Co => 
                           q_1_1_42_port);
   HA_L_0_0_42 : HA_42 port map( A => X_Logic1_port, B => q_0_1_42_port, S => 
                           q_1_0_42_port, C => q_1_0_43_port);
   HA_R_0_3_26 : HA_41 port map( A => q_0_3_26_port, B => q_0_4_26_port, S => 
                           q_1_2_26_port, C => q_1_3_27_port);
   HA_R_0_3_27 : HA_40 port map( A => q_0_3_27_port, B => q_0_4_27_port, S => 
                           n357, C => q_1_3_28_port);
   FA_C_0_3_28 : FA_592 port map( A => q_0_3_28_port, B => q_0_4_28_port, Ci =>
                           q_0_5_28_port, S => q_1_2_28_port, Co => n347);
   FA_C_0_3_29 : FA_591 port map( A => q_0_3_29_port, B => q_0_4_29_port, Ci =>
                           q_0_5_29_port, S => q_1_2_29_port, Co => 
                           q_1_3_30_port);
   FA_C_0_3_30 : FA_590 port map( A => q_0_3_30_port, B => q_0_4_30_port, Ci =>
                           q_0_5_30_port, S => q_1_2_30_port, Co => 
                           q_1_3_31_port);
   FA_C_0_3_31 : FA_589 port map( A => q_0_3_31_port, B => q_0_4_31_port, Ci =>
                           q_0_5_31_port, S => q_1_2_31_port, Co => 
                           q_1_3_32_port);
   FA_C_0_3_32 : FA_588 port map( A => q_0_3_32_port, B => q_0_4_32_port, Ci =>
                           q_0_5_32_port, S => q_1_2_32_port, Co => 
                           q_1_3_33_port);
   FA_C_0_3_33 : FA_587 port map( A => q_0_3_33_port, B => q_0_4_33_port, Ci =>
                           q_0_5_33_port, S => q_1_2_33_port, Co => 
                           q_1_3_34_port);
   FA_C_0_3_34 : FA_586 port map( A => q_0_3_34_port, B => q_0_4_34_port, Ci =>
                           q_0_5_34_port, S => q_1_2_34_port, Co => 
                           q_1_3_35_port);
   FA_C_0_3_35 : FA_585 port map( A => q_0_3_35_port, B => q_0_4_35_port, Ci =>
                           q_0_5_35_port, S => q_1_2_35_port, Co => 
                           q_1_3_36_port);
   FA_C_0_3_36 : FA_584 port map( A => q_0_3_36_port, B => q_0_4_36_port, Ci =>
                           q_0_5_36_port, S => q_1_2_36_port, Co => 
                           q_1_3_37_port);
   FA_C_0_3_37 : FA_583 port map( A => q_0_3_37_port, B => q_0_4_37_port, Ci =>
                           q_0_5_37_port, S => q_1_2_37_port, Co => 
                           q_1_3_38_port);
   FA_C_0_3_38 : FA_582 port map( A => q_0_3_38_port, B => q_0_4_38_port, Ci =>
                           q_0_5_38_port, S => q_1_2_38_port, Co => 
                           q_1_3_39_port);
   FA_C_0_3_39 : FA_581 port map( A => q_0_3_39_port, B => q_0_4_39_port, Ci =>
                           q_0_5_39_port, S => q_1_2_39_port, Co => 
                           q_1_3_40_port);
   HA_L_0_3_40 : HA_39 port map( A => q_0_3_40_port, B => q_0_4_40_port, S => 
                           q_1_2_40_port, C => q_1_2_41_port);
   HA_R_0_6_28 : HA_38 port map( A => q_0_6_28_port, B => q_0_7_28_port, S => 
                           q_1_4_28_port, C => q_1_5_29_port);
   HA_R_0_6_29 : HA_37 port map( A => q_0_6_29_port, B => q_0_7_29_port, S => 
                           q_1_4_29_port, C => q_1_5_30_port);
   FA_C_0_6_30 : FA_580 port map( A => q_0_6_30_port, B => q_0_7_30_port, Ci =>
                           q_0_8_30_port, S => q_1_4_30_port, Co => 
                           q_1_5_31_port);
   FA_C_0_6_31 : FA_579 port map( A => q_0_6_31_port, B => q_0_7_31_port, Ci =>
                           q_0_8_31_port, S => q_1_4_31_port, Co => 
                           q_1_5_32_port);
   FA_C_0_6_32 : FA_578 port map( A => q_0_6_32_port, B => q_0_7_32_port, Ci =>
                           q_0_8_32_port, S => q_1_4_32_port, Co => 
                           q_1_5_33_port);
   FA_C_0_6_33 : FA_577 port map( A => q_0_6_33_port, B => q_0_7_33_port, Ci =>
                           q_0_8_33_port, S => q_1_4_33_port, Co => 
                           q_1_5_34_port);
   FA_C_0_6_34 : FA_576 port map( A => q_0_6_34_port, B => q_0_7_34_port, Ci =>
                           q_0_8_34_port, S => q_1_4_34_port, Co => 
                           q_1_5_35_port);
   FA_C_0_6_35 : FA_575 port map( A => q_0_6_35_port, B => q_0_7_35_port, Ci =>
                           q_0_8_35_port, S => q_1_4_35_port, Co => 
                           q_1_5_36_port);
   FA_C_0_6_36 : FA_574 port map( A => q_0_6_36_port, B => q_0_7_36_port, Ci =>
                           q_0_8_36_port, S => q_1_4_36_port, Co => 
                           q_1_5_37_port);
   FA_C_0_6_37 : FA_573 port map( A => q_0_6_37_port, B => q_0_7_37_port, Ci =>
                           q_0_8_37_port, S => q_1_4_37_port, Co => 
                           q_1_5_38_port);
   HA_L_0_6_38 : HA_36 port map( A => q_0_6_38_port, B => q_0_7_38_port, S => 
                           q_1_4_38_port, C => q_1_4_39_port);
   HA_R_0_9_30 : HA_35 port map( A => q_0_9_30_port, B => q_0_10_30_port, S => 
                           q_1_6_30_port, C => q_1_7_31_port);
   HA_R_0_9_31 : HA_34 port map( A => q_0_9_31_port, B => q_0_10_31_port, S => 
                           q_1_6_31_port, C => q_1_7_32_port);
   FA_C_0_9_32 : FA_572 port map( A => q_0_9_32_port, B => q_0_10_32_port, Ci 
                           => q_0_11_32_port, S => q_1_6_32_port, Co => 
                           q_1_7_33_port);
   FA_C_0_9_33 : FA_571 port map( A => q_0_9_33_port, B => q_0_10_33_port, Ci 
                           => q_0_11_33_port, S => q_1_6_33_port, Co => 
                           q_1_7_34_port);
   FA_C_0_9_34 : FA_570 port map( A => q_0_9_34_port, B => q_0_10_34_port, Ci 
                           => q_0_11_34_port, S => q_1_6_34_port, Co => 
                           q_1_7_35_port);
   FA_C_0_9_35 : FA_569 port map( A => q_0_9_35_port, B => q_0_10_35_port, Ci 
                           => q_0_11_35_port, S => q_1_6_35_port, Co => 
                           q_1_7_36_port);
   HA_L_0_9_36 : HA_33 port map( A => q_0_9_36_port, B => q_0_10_36_port, S => 
                           q_1_6_36_port, C => q_1_6_37_port);
   HA_R_1_0_16 : HA_32 port map( A => q_0_0_16_port, B => q_0_1_16_port, S => 
                           q_2_0_16_port, C => q_2_1_17_port);
   HA_R_1_0_17 : HA_31 port map( A => q_0_0_17_port, B => q_0_1_17_port, S => 
                           q_2_0_17_port, C => q_2_1_18_port);
   FA_C_1_0_18 : FA_568 port map( A => q_0_0_18_port, B => q_0_1_18_port, Ci =>
                           q_0_2_18_port, S => q_2_0_18_port, Co => 
                           q_2_1_19_port);
   FA_C_1_0_19 : FA_567 port map( A => q_0_0_19_port, B => q_0_1_19_port, Ci =>
                           q_0_2_19_port, S => q_2_0_19_port, Co => 
                           q_2_1_20_port);
   FA_C_1_0_20 : FA_566 port map( A => q_0_0_20_port, B => q_0_1_20_port, Ci =>
                           q_0_2_20_port, S => q_2_0_20_port, Co => 
                           q_2_1_21_port);
   FA_C_1_0_21 : FA_565 port map( A => q_0_0_21_port, B => q_0_1_21_port, Ci =>
                           q_0_2_21_port, S => q_2_0_21_port, Co => 
                           q_2_1_22_port);
   FA_C_1_0_22 : FA_564 port map( A => q_0_0_22_port, B => n362, Ci => 
                           q_0_2_22_port, S => q_2_0_22_port, Co => 
                           q_2_1_23_port);
   FA_C_1_0_23 : FA_563 port map( A => q_0_0_23_port, B => q_0_1_23_port, Ci =>
                           q_0_2_23_port, S => q_2_0_23_port, Co => 
                           q_2_1_24_port);
   FA_C_1_0_24 : FA_562 port map( A => q_1_0_24_port, B => q_0_2_24_port, Ci =>
                           q_0_3_24_port, S => q_2_0_24_port, Co => 
                           q_2_1_25_port);
   FA_C_1_0_25 : FA_561 port map( A => q_1_0_25_port, B => q_1_1_25_port, Ci =>
                           q_0_2_25_port, S => q_2_0_25_port, Co => 
                           q_2_1_26_port);
   FA_C_1_0_26 : FA_560 port map( A => q_1_0_26_port, B => q_1_1_26_port, Ci =>
                           q_1_2_26_port, S => q_2_0_26_port, Co => 
                           q_2_1_27_port);
   FA_C_1_0_27 : FA_559 port map( A => q_1_0_27_port, B => n351, Ci => n357, S 
                           => q_2_0_27_port, Co => q_2_1_28_port, clk => clk);
   FA_C_1_0_28 : FA_558 port map( A => n348, B => q_1_1_28_port, Ci => 
                           q_1_2_28_port, S => q_2_0_28_port, Co => 
                           q_2_1_29_port);
   FA_C_1_0_29 : FA_557 port map( A => n352, B => q_1_1_29_port, Ci => 
                           q_1_2_29_port, S => q_2_0_29_port, Co => 
                           q_2_1_30_port);
   FA_C_1_0_30 : FA_556 port map( A => q_1_0_30_port, B => q_1_1_30_port, Ci =>
                           q_1_2_30_port, S => q_2_0_30_port, Co => 
                           q_2_1_31_port);
   FA_C_1_0_31 : FA_555 port map( A => q_1_0_31_port, B => q_1_1_31_port, Ci =>
                           q_1_2_31_port, S => q_2_0_31_port, Co => 
                           q_2_1_32_port, clk => clk);
   FA_C_1_0_32 : FA_554 port map( A => q_1_0_32_port, B => q_1_1_32_port, Ci =>
                           q_1_2_32_port, S => q_2_0_32_port, Co => 
                           q_2_1_33_port, clk => clk);
   FA_C_1_0_33 : FA_553 port map( A => q_1_0_33_port, B => q_1_1_33_port, Ci =>
                           q_1_2_33_port, S => q_2_0_33_port, Co => 
                           q_2_1_34_port, clk => clk);
   FA_C_1_0_34 : FA_552 port map( A => q_1_0_34_port, B => q_1_1_34_port, Ci =>
                           q_1_2_34_port, S => n374, Co => q_2_1_35_port, clk 
                           => clk);
   FA_C_1_0_35 : FA_551 port map( A => q_1_0_35_port, B => q_1_1_35_port, Ci =>
                           q_1_2_35_port, S => q_2_0_35_port, Co => 
                           q_2_1_36_port, clk => clk);
   FA_C_1_0_36 : FA_550 port map( A => q_1_0_36_port, B => q_1_1_36_port, Ci =>
                           q_1_2_36_port, S => q_2_0_36_port, Co => 
                           q_2_1_37_port);
   FA_C_1_0_37 : FA_549 port map( A => q_1_0_37_port, B => q_1_1_37_port, Ci =>
                           q_1_2_37_port, S => q_2_0_37_port, Co => 
                           q_2_1_38_port, clk => clk);
   FA_C_1_0_38 : FA_548 port map( A => q_1_0_38_port, B => q_1_1_38_port, Ci =>
                           q_1_2_38_port, S => q_2_0_38_port, Co => 
                           q_2_1_39_port, clk => clk);
   FA_C_1_0_39 : FA_547 port map( A => q_1_0_39_port, B => q_1_1_39_port, Ci =>
                           q_1_2_39_port, S => q_2_0_39_port, Co => 
                           q_2_1_40_port, clk => clk);
   FA_C_1_0_40 : FA_546 port map( A => q_1_0_40_port, B => q_1_1_40_port, Ci =>
                           q_1_2_40_port, S => n377, Co => q_2_1_41_port, clk 
                           => clk);
   FA_C_1_0_41 : FA_545 port map( A => q_1_0_41_port, B => q_1_1_41_port, Ci =>
                           q_1_2_41_port, S => q_2_0_41_port, Co => 
                           q_2_1_42_port);
   FA_C_1_0_42 : FA_544 port map( A => q_1_0_42_port, B => q_1_1_42_port, Ci =>
                           q_0_2_42_port, S => q_2_0_42_port, Co => 
                           q_2_1_43_port);
   FA_C_1_0_43 : FA_543 port map( A => q_1_0_43_port, Ci => q_0_1_43_port, S =>
                           q_2_0_43_port, Co => q_2_1_44_port, B_BAR => B(11));
   FA_C_1_0_44 : FA_542 port map( A => X_Logic1_port, B => q_0_1_44_port, Ci =>
                           q_0_2_44_port, S => q_2_0_44_port, Co => 
                           q_2_1_45_port);
   FA_C_1_0_45 : FA_541 port map( B => q_0_1_45_port, Ci => q_0_2_45_port, S =>
                           q_2_0_45_port, Co => q_2_1_46_port, A_BAR => B(13));
   FA_C_1_0_46 : FA_540 port map( A => X_Logic1_port, B => q_0_1_46_port, Ci =>
                           q_0_2_46_port, S => q_2_0_46_port, Co => 
                           q_2_1_47_port);
   FA_C_1_0_47 : FA_539 port map( B => q_0_1_47_port, Ci => q_0_2_47_port, S =>
                           q_2_0_47_port, Co => n_2032, A => B(15));
   HA_R_1_3_18 : HA_29 port map( A => q_0_3_18_port, B => q_0_4_18_port, S => 
                           q_2_2_18_port, C => q_2_3_19_port);
   HA_R_1_3_19 : HA_28 port map( A => q_0_3_19_port, B => q_0_4_19_port, S => 
                           q_2_2_19_port, C => q_2_3_20_port);
   FA_C_1_3_20 : FA_536 port map( A => q_0_3_20_port, B => q_0_4_20_port, Ci =>
                           q_0_5_20_port, S => q_2_2_20_port, Co => 
                           q_2_3_21_port);
   FA_C_1_3_21 : FA_535 port map( A => q_0_3_21_port, B => q_0_4_21_port, Ci =>
                           q_0_5_21_port, S => q_2_2_21_port, Co => 
                           q_2_3_22_port);
   FA_C_1_3_22 : FA_534 port map( A => q_0_3_22_port, B => q_0_4_22_port, Ci =>
                           q_0_5_22_port, S => q_2_2_22_port, Co => 
                           q_2_3_23_port);
   FA_C_1_3_23 : FA_533 port map( A => q_0_3_23_port, B => q_0_4_23_port, Ci =>
                           q_0_5_23_port, S => q_2_2_23_port, Co => 
                           q_2_3_24_port);
   FA_C_1_3_24 : FA_532 port map( A => q_0_4_24_port, B => q_0_5_24_port, Ci =>
                           q_0_6_24_port, S => q_2_2_24_port, Co => 
                           q_2_3_25_port);
   FA_C_1_3_25 : FA_531 port map( A => q_0_3_25_port, B => q_0_4_25_port, Ci =>
                           q_0_5_25_port, S => q_2_2_25_port, Co => 
                           q_2_3_26_port);
   FA_C_1_3_26 : FA_530 port map( A => q_0_5_26_port, B => q_0_6_26_port, Ci =>
                           q_0_7_26_port, S => q_2_2_26_port, Co => 
                           q_2_3_27_port, clk => clk);
   FA_C_1_3_27 : FA_529 port map( A => q_1_3_27_port, B => q_0_5_27_port, Ci =>
                           q_0_6_27_port, S => q_2_2_27_port, Co => 
                           q_2_3_28_port);
   FA_C_1_3_28 : FA_528 port map( A => q_1_3_28_port, B => q_1_4_28_port, Ci =>
                           q_0_8_28_port, S => q_2_2_28_port, Co => 
                           q_2_3_29_port);
   FA_C_1_3_29 : FA_527 port map( A => n347, B => q_1_4_29_port, Ci => 
                           q_1_5_29_port, S => q_2_2_29_port, Co => 
                           q_2_3_30_port);
   FA_C_1_3_30 : FA_526 port map( A => q_1_3_30_port, B => q_1_4_30_port, Ci =>
                           q_1_5_30_port, S => q_2_2_30_port, Co => 
                           q_2_3_31_port, clk => clk);
   FA_C_1_3_31 : FA_525 port map( A => q_1_3_31_port, B => q_1_4_31_port, Ci =>
                           q_1_5_31_port, S => q_2_2_31_port, Co => 
                           q_2_3_32_port, clk => clk);
   FA_C_1_3_32 : FA_524 port map( A => q_1_3_32_port, B => q_1_4_32_port, S => 
                           q_2_2_32_port, Co => n365, clk => clk, Ci_BAR => 
                           q_1_5_32_port);
   FA_C_1_3_33 : FA_523 port map( A => q_1_3_33_port, B => q_1_4_33_port, Ci =>
                           q_1_5_33_port, S => q_2_2_33_port, Co => 
                           q_2_3_34_port, clk => clk);
   FA_C_1_3_34 : FA_522 port map( A => q_1_3_34_port, B => q_1_4_34_port, Ci =>
                           q_1_5_34_port, S => q_2_2_34_port, Co => 
                           q_2_3_35_port, clk => clk);
   FA_C_1_3_35 : FA_521 port map( A => q_1_3_35_port, B => q_1_4_35_port, Ci =>
                           q_1_5_35_port, S => q_2_2_35_port, Co => 
                           q_2_3_36_port, clk => clk);
   FA_C_1_3_36 : FA_520 port map( A => q_1_3_36_port, B => q_1_4_36_port, Ci =>
                           q_1_5_36_port, S => q_2_2_36_port, Co => 
                           q_2_3_37_port, clk => clk);
   FA_C_1_3_37 : FA_519 port map( A => q_1_3_37_port, B => q_1_4_37_port, Ci =>
                           q_1_5_37_port, S => q_2_2_37_port, Co => 
                           q_2_3_38_port, clk => clk);
   FA_C_1_3_38 : FA_518 port map( A => q_1_3_38_port, B => q_1_4_38_port, Ci =>
                           q_1_5_38_port, S => n363, Co => q_2_3_39_port, clk 
                           => clk);
   FA_C_1_3_39 : FA_517 port map( A => q_1_3_39_port, B => q_1_4_39_port, Ci =>
                           q_0_6_39_port, S => q_2_2_39_port, Co => 
                           q_2_3_40_port);
   FA_C_1_3_40 : FA_516 port map( A => q_1_3_40_port, B => q_0_5_40_port, Ci =>
                           q_0_6_40_port, S => q_2_2_40_port, Co => 
                           q_2_3_41_port, clk => clk);
   FA_C_1_3_41 : FA_515 port map( A => q_0_3_41_port, B => q_0_4_41_port, Ci =>
                           q_0_5_41_port, S => q_2_2_41_port, Co => 
                           q_2_3_42_port);
   FA_C_1_3_42 : FA_514 port map( A => q_0_3_42_port, B => q_0_4_42_port, Ci =>
                           q_0_5_42_port, S => q_2_2_42_port, Co => 
                           q_2_3_43_port);
   FA_C_1_3_43 : FA_513 port map( A => q_0_2_43_port, B => q_0_3_43_port, Ci =>
                           q_0_4_43_port, S => q_2_2_43_port, Co => 
                           q_2_3_44_port);
   FA_C_1_3_44 : FA_512 port map( A => q_0_3_44_port, B => q_0_4_44_port, Ci =>
                           q_0_5_44_port, S => q_2_2_44_port, Co => 
                           q_2_3_45_port);
   FA_C_1_3_45 : FA_511 port map( A => q_0_3_45_port, B => q_0_4_45_port, Ci =>
                           q_0_5_45_port, S => q_2_2_45_port, Co => 
                           q_2_3_46_port);
   FA_C_1_3_46 : FA_510 port map( A => q_0_3_46_port, B => q_0_4_46_port, Ci =>
                           q_0_5_46_port, S => q_2_2_46_port, Co => 
                           q_2_3_47_port);
   FA_C_1_3_47 : FA_509 port map( A => q_0_3_47_port, B => q_0_4_47_port, Ci =>
                           q_0_5_47_port, S => q_2_2_47_port, Co => n_2033);
   HA_R_1_6_20 : HA_26 port map( A => q_0_6_20_port, B => q_0_7_20_port, S => 
                           q_2_4_20_port, C => q_2_5_21_port);
   HA_R_1_6_21 : HA_25 port map( A => q_0_6_21_port, B => q_0_7_21_port, S => 
                           q_2_4_21_port, C => q_2_5_22_port);
   FA_C_1_6_22 : FA_508 port map( A => q_0_6_22_port, B => q_0_7_22_port, Ci =>
                           q_0_8_22_port, S => q_2_4_22_port, Co => 
                           q_2_5_23_port);
   FA_C_1_6_23 : FA_507 port map( A => q_0_6_23_port, B => q_0_7_23_port, Ci =>
                           q_0_8_23_port, S => q_2_4_23_port, Co => 
                           q_2_5_24_port);
   FA_C_1_6_24 : FA_506 port map( A => q_0_7_24_port, B => q_0_8_24_port, Ci =>
                           q_0_9_24_port, S => q_2_4_24_port, Co => 
                           q_2_5_25_port);
   FA_C_1_6_25 : FA_505 port map( A => q_0_6_25_port, B => q_0_7_25_port, Ci =>
                           q_0_8_25_port, S => q_2_4_25_port, Co => 
                           q_2_5_26_port);
   FA_C_1_6_26 : FA_504 port map( A => q_0_8_26_port, B => q_0_9_26_port, Ci =>
                           q_0_10_26_port, S => q_2_4_26_port, Co => 
                           q_2_5_27_port);
   FA_C_1_6_27 : FA_503 port map( A => q_0_7_27_port, B => q_0_8_27_port, Ci =>
                           q_0_9_27_port, S => q_2_4_27_port, Co => 
                           q_2_5_28_port);
   FA_C_1_6_28 : FA_502 port map( A => q_0_9_28_port, B => q_0_10_28_port, Ci 
                           => q_0_11_28_port, S => q_2_4_28_port, Co => 
                           q_2_5_29_port);
   FA_C_1_6_29 : FA_501 port map( A => q_0_8_29_port, B => n361, Ci => 
                           q_0_10_29_port, S => q_2_4_29_port, Co => 
                           q_2_5_30_port);
   FA_C_1_6_30 : FA_500 port map( A => q_1_6_30_port, B => q_0_11_30_port, Ci 
                           => q_0_12_30_port, S => q_2_4_30_port, Co => 
                           q_2_5_31_port);
   FA_C_1_6_31 : FA_499 port map( A => q_1_6_31_port, B => q_1_7_31_port, Ci =>
                           q_0_11_31_port, S => q_2_4_31_port, Co => 
                           q_2_5_32_port);
   FA_C_1_6_32 : FA_498 port map( A => q_1_6_32_port, B => q_1_7_32_port, Ci =>
                           q_0_12_32_port, S => q_2_4_32_port, Co => 
                           q_2_5_33_port);
   FA_C_1_6_33 : FA_497 port map( A => q_1_6_33_port, B => q_1_7_33_port, Ci =>
                           q_0_12_33_port, S => q_2_4_33_port, Co => 
                           q_2_5_34_port, clk => clk);
   FA_C_1_6_34 : FA_496 port map( A => q_1_6_34_port, B => q_1_7_34_port, Ci =>
                           q_0_12_34_port, S => q_2_4_34_port, Co => 
                           q_2_5_35_port);
   FA_C_1_6_35 : FA_495 port map( A => q_1_6_35_port, B => q_1_7_35_port, Ci =>
                           q_0_12_35_port, S => q_2_4_35_port, Co => 
                           q_2_5_36_port, clk => clk);
   FA_C_1_6_36 : FA_494 port map( A => q_1_6_36_port, B => q_1_7_36_port, Ci =>
                           q_0_11_36_port, S => q_2_4_36_port, Co => 
                           q_2_5_37_port);
   FA_C_1_6_37 : FA_493 port map( A => q_1_6_37_port, B => q_0_9_37_port, S => 
                           q_2_4_37_port, Co => q_2_5_38_port, Ci_BAR => 
                           q_0_10_37_port);
   FA_C_1_6_38 : FA_492 port map( A => q_0_8_38_port, B => q_0_9_38_port, S => 
                           q_2_4_38_port, Co => q_2_5_39_port, Ci_BAR => 
                           q_0_10_38_port);
   FA_C_1_6_39 : FA_491 port map( A => q_0_7_39_port, B => q_0_8_39_port, S => 
                           q_2_4_39_port, Co => q_2_5_40_port, Ci_BAR => 
                           q_0_9_39_port);
   FA_C_1_6_40 : FA_490 port map( A => q_0_7_40_port, B => q_0_8_40_port, S => 
                           q_2_4_40_port, Co => q_2_5_41_port, Ci_BAR => 
                           q_0_9_40_port);
   FA_C_1_6_41 : FA_489 port map( A => q_0_6_41_port, B => q_0_7_41_port, S => 
                           q_2_4_41_port, Co => q_2_5_42_port, Ci_BAR => 
                           q_0_8_41_port);
   FA_C_1_6_42 : FA_488 port map( A => q_0_6_42_port, B => q_0_7_42_port, S => 
                           q_2_4_42_port, Co => q_2_5_43_port, Ci_BAR => 
                           q_0_8_42_port);
   FA_C_1_6_43 : FA_487 port map( A => q_0_5_43_port, B => q_0_6_43_port, S => 
                           q_2_4_43_port, Co => q_2_5_44_port, Ci_BAR => 
                           q_0_7_43_port);
   FA_C_1_6_44 : FA_486 port map( A => q_0_6_44_port, Ci => net102806, Co => 
                           q_2_5_45_port, B_BAR => q_0_7_44_port, S_BAR => 
                           q_2_4_44_port);
   FA_C_1_6_45 : FA_485 port map( B => net102804, Ci => net102805, Co => n_2034
                           , A_BAR => q_0_6_45_port, S_BAR => q_2_4_45_port);
   HA_L_1_6_46 : HA_24 port map( B => net102803, C => n_2035, S_BAR => 
                           q_2_4_46_port, A_BAR => q_0_6_46_port);
   HA_R_1_9_22 : HA_23 port map( A => q_0_9_22_port, B => q_0_10_22_port, S => 
                           q_2_6_22_port, C => q_2_7_23_port);
   HA_R_1_9_23 : HA_22 port map( A => q_0_9_23_port, B => q_0_10_23_port, S => 
                           n356, C => q_2_7_24_port);
   FA_C_1_9_24 : FA_484 port map( A => q_0_10_24_port, B => q_0_11_24_port, Ci 
                           => q_0_12_24_port, S => q_2_6_24_port, Co => 
                           q_2_7_25_port);
   FA_C_1_9_25 : FA_483 port map( A => q_0_9_25_port, B => q_0_10_25_port, Ci 
                           => q_0_11_25_port, S => q_2_6_25_port, Co => 
                           q_2_7_26_port);
   FA_C_1_9_26 : FA_482 port map( A => q_0_11_26_port, Ci => net102802, S => 
                           q_2_6_26_port, Co => q_2_7_27_port, B_BAR => 
                           q_0_12_26_port);
   FA_C_1_9_27 : FA_481 port map( A => q_0_10_27_port, B => q_0_11_27_port, Ci 
                           => q_0_12_27_port, S => q_2_6_27_port, Co => 
                           q_2_7_28_port);
   FA_C_1_9_28 : FA_480 port map( B => net102800, Ci => net102801, S => 
                           q_2_6_28_port, Co => n_2036, A_BAR => q_0_12_28_port
                           );
   FA_C_1_9_29 : FA_479 port map( A => q_0_11_29_port, Ci => net102799, S => 
                           q_2_6_29_port, Co => q_2_7_30_port, B_BAR => 
                           q_0_12_29_port);
   FA_C_1_9_31 : FA_477 port map( B => net102797, Ci => net102798, Co => n_2037
                           , A_BAR => q_0_12_31_port, S_BAR => q_2_6_31_port);
   HA_R_2_0_10 : HA_20 port map( A => q_0_0_10_port, B => q_0_1_10_port, S => 
                           n355, C => q_3_1_11_port);
   HA_R_2_0_11 : HA_19 port map( A => q_0_0_11_port, B => q_0_1_11_port, S => 
                           n354, C => q_3_1_12_port);
   FA_C_2_0_12 : FA_464 port map( A => q_0_0_12_port, B => q_0_1_12_port, Ci =>
                           q_0_2_12_port, S => q_3_0_12_port, Co => 
                           q_3_1_13_port);
   FA_C_2_0_13 : FA_463 port map( A => q_0_0_13_port, B => q_0_1_13_port, Ci =>
                           q_0_2_13_port, S => q_3_0_13_port, Co => 
                           q_3_1_14_port);
   FA_C_2_0_14 : FA_462 port map( A => q_0_0_14_port, B => q_0_1_14_port, Ci =>
                           q_0_2_14_port, S => q_3_0_14_port, Co => 
                           q_3_1_15_port);
   FA_C_2_0_15 : FA_461 port map( A => q_0_0_15_port, B => q_0_1_15_port, Ci =>
                           q_0_2_15_port, S => q_3_0_15_port, Co => 
                           q_3_1_16_port);
   FA_C_2_0_16 : FA_460 port map( A => q_2_0_16_port, B => q_0_2_16_port, Ci =>
                           q_0_3_16_port, S => q_3_0_16_port, Co => 
                           q_3_1_17_port);
   FA_C_2_0_17 : FA_459 port map( A => q_2_0_17_port, B => q_2_1_17_port, Ci =>
                           q_0_2_17_port, S => q_3_0_17_port, Co => 
                           q_3_1_18_port, clk => clk);
   FA_C_2_0_18 : FA_458 port map( A => q_2_0_18_port, B => q_2_1_18_port, Ci =>
                           q_2_2_18_port, S => q_3_0_18_port, Co => 
                           q_3_1_19_port, clk => clk);
   FA_C_2_0_19 : FA_457 port map( A => q_2_0_19_port, B => q_2_1_19_port, Ci =>
                           q_2_2_19_port, S => q_3_0_19_port, Co => 
                           q_3_1_20_port, clk => clk);
   FA_C_2_0_20 : FA_456 port map( A => q_2_0_20_port, B => q_2_1_20_port, Ci =>
                           q_2_2_20_port, S => q_3_0_20_port, Co => 
                           q_3_1_21_port, clk => clk);
   FA_C_2_0_21 : FA_455 port map( A => q_2_0_21_port, B => q_2_1_21_port, Ci =>
                           q_2_2_21_port, S => q_3_0_21_port, Co => 
                           q_3_1_22_port, clk => clk);
   FA_C_2_0_22 : FA_454 port map( A => q_2_0_22_port, B => q_2_1_22_port, Ci =>
                           q_2_2_22_port, S => q_3_0_22_port, Co => 
                           q_3_1_23_port, clk => clk);
   FA_C_2_0_23 : FA_453 port map( A => q_2_0_23_port, B => q_2_1_23_port, Ci =>
                           q_2_2_23_port, S => n373, Co => q_3_1_24_port, clk 
                           => clk);
   FA_C_2_0_24 : FA_452 port map( A => q_2_0_24_port, B => q_2_1_24_port, Ci =>
                           q_2_2_24_port, S => q_3_0_24_port, Co => 
                           q_3_1_25_port, clk => clk);
   FA_C_2_0_25 : FA_451 port map( A => q_2_0_25_port, B => q_2_1_25_port, Ci =>
                           q_2_2_25_port, S => q_3_0_25_port, Co => 
                           q_3_1_26_port, clk => clk);
   FA_C_2_0_26 : FA_450 port map( A => q_2_0_26_port, B => q_2_1_26_port, Ci =>
                           q_2_2_26_port, S => q_3_0_26_port, Co => 
                           q_3_1_27_port, clk => clk);
   FA_C_2_0_27 : FA_449 port map( A => q_2_0_27_port, B => q_2_1_27_port, Ci =>
                           q_2_2_27_port, S => q_3_0_27_port, Co => 
                           q_3_1_28_port, clk => clk);
   FA_C_2_0_28 : FA_448 port map( A => q_2_0_28_port, B => q_2_1_28_port, Ci =>
                           q_2_2_28_port, S => q_3_0_28_port, Co => 
                           q_3_1_29_port, clk => clk);
   FA_C_2_0_29 : FA_447 port map( A => q_2_0_29_port, B => q_2_1_29_port, Ci =>
                           q_2_2_29_port, S => q_3_0_29_port, Co => 
                           q_3_1_30_port, clk => clk);
   FA_C_2_0_30 : FA_446 port map( A => q_2_0_30_port, B => q_2_1_30_port, Ci =>
                           q_2_2_30_port, S => q_3_0_30_port, Co => 
                           q_3_1_31_port, clk => clk);
   FA_C_2_0_31 : FA_445 port map( A => q_2_0_31_port, B => q_2_1_31_port, Ci =>
                           q_2_2_31_port, S => q_3_0_31_port, Co => 
                           q_3_1_32_port, clk => clk);
   FA_C_2_0_32 : FA_444 port map( A => q_2_0_32_port, B => q_2_1_32_port, Ci =>
                           q_2_2_32_port, S => q_3_0_32_port, Co => 
                           q_3_1_33_port);
   FA_C_2_0_33 : FA_443 port map( A => q_2_0_33_port, B => q_2_1_33_port, Ci =>
                           q_2_2_33_port, S => q_3_0_33_port, Co => 
                           q_3_1_34_port, clk => clk);
   FA_C_2_0_34 : FA_442 port map( A => n374, B => q_2_1_34_port, Ci => 
                           q_2_2_34_port, S => q_3_0_34_port, Co => n353);
   FA_C_2_0_35 : FA_441 port map( A => q_2_0_35_port, B => q_2_1_35_port, Ci =>
                           q_2_2_35_port, S => q_3_0_35_port, Co => 
                           q_3_1_36_port, clk => clk);
   FA_C_2_0_36 : FA_440 port map( A => q_2_0_36_port, B => q_2_1_36_port, Ci =>
                           q_2_2_36_port, S => q_3_0_36_port, Co => 
                           q_3_1_37_port, clk => clk);
   FA_C_2_0_37 : FA_439 port map( A => q_2_0_37_port, B => q_2_1_37_port, Ci =>
                           q_2_2_37_port, S => q_3_0_37_port, Co => 
                           q_3_1_38_port, clk => clk);
   FA_C_2_0_38 : FA_438 port map( A => q_2_0_38_port, B => q_2_1_38_port, Ci =>
                           n363, S => q_3_0_38_port, Co => q_3_1_39_port);
   FA_C_2_0_39 : FA_437 port map( A => q_2_0_39_port, B => q_2_1_39_port, Ci =>
                           q_2_2_39_port, S => q_3_0_39_port, Co => 
                           q_3_1_40_port, clk => clk);
   FA_C_2_0_40 : FA_436 port map( A => n377, B => q_2_1_40_port, Ci => 
                           q_2_2_40_port, S => q_3_0_40_port, Co => 
                           q_3_1_41_port);
   FA_C_2_0_41 : FA_435 port map( A => q_2_0_41_port, B => q_2_1_41_port, Ci =>
                           q_2_2_41_port, S => q_3_0_41_port, Co => 
                           q_3_1_42_port, clk => clk);
   FA_C_2_0_42 : FA_434 port map( A => q_2_0_42_port, B => q_2_1_42_port, Ci =>
                           q_2_2_42_port, S => q_3_0_42_port, Co => 
                           q_3_1_43_port, clk => clk);
   FA_C_2_0_43 : FA_433 port map( A => q_2_0_43_port, B => q_2_1_43_port, Ci =>
                           q_2_2_43_port, S => n367, Co => n368, clk => clk);
   FA_C_2_0_44 : FA_432 port map( A => q_2_0_44_port, B => q_2_1_44_port, Ci =>
                           q_2_2_44_port, S => q_3_0_44_port, Co => 
                           q_3_1_45_port, clk => clk);
   FA_C_2_0_45 : FA_431 port map( A => q_2_0_45_port, B => q_2_1_45_port, Ci =>
                           q_2_2_45_port, S => q_3_0_45_port, Co => 
                           q_3_1_46_port, clk => clk);
   FA_C_2_0_46 : FA_430 port map( A => q_2_0_46_port, B => q_2_1_46_port, Ci =>
                           q_2_2_46_port, S => q_3_0_46_port, Co => 
                           q_3_1_47_port, clk => clk);
   FA_C_2_0_47 : FA_429 port map( A => q_2_0_47_port, B => q_2_1_47_port, Ci =>
                           q_2_2_47_port, S => q_3_0_47_port, Co => n_2038, clk
                           => clk);
   HA_R_2_3_12 : HA_17 port map( A => q_0_3_12_port, B => q_0_4_12_port, S => 
                           q_3_2_12_port, C => q_3_3_13_port);
   HA_R_2_3_13 : HA_16 port map( A => q_0_3_13_port, B => q_0_4_13_port, S => 
                           q_3_2_13_port, C => q_3_3_14_port);
   FA_C_2_3_14 : FA_420 port map( A => q_0_3_14_port, B => q_0_4_14_port, Ci =>
                           q_0_5_14_port, S => q_3_2_14_port, Co => 
                           q_3_3_15_port);
   FA_C_2_3_15 : FA_419 port map( A => q_0_3_15_port, B => q_0_4_15_port, Ci =>
                           q_0_5_15_port, S => q_3_2_15_port, Co => 
                           q_3_3_16_port);
   FA_C_2_3_16 : FA_418 port map( A => q_0_4_16_port, B => q_0_5_16_port, Ci =>
                           q_0_6_16_port, S => q_3_2_16_port, Co => 
                           q_3_3_17_port);
   FA_C_2_3_17 : FA_417 port map( A => q_0_3_17_port, B => q_0_4_17_port, Ci =>
                           q_0_5_17_port, S => q_3_2_17_port, Co => 
                           q_3_3_18_port);
   FA_C_2_3_18 : FA_416 port map( A => q_0_5_18_port, B => q_0_6_18_port, Ci =>
                           q_0_7_18_port, S => q_3_2_18_port, Co => 
                           q_3_3_19_port);
   FA_C_2_3_19 : FA_415 port map( A => q_2_3_19_port, B => q_0_5_19_port, Ci =>
                           q_0_6_19_port, S => q_3_2_19_port, Co => 
                           q_3_3_20_port);
   FA_C_2_3_20 : FA_414 port map( A => q_2_3_20_port, B => q_2_4_20_port, Ci =>
                           q_0_8_20_port, S => q_3_2_20_port, Co => 
                           q_3_3_21_port, clk => clk);
   FA_C_2_3_21 : FA_413 port map( A => q_2_3_21_port, B => q_2_4_21_port, Ci =>
                           q_2_5_21_port, S => n370, Co => q_3_3_22_port, clk 
                           => clk);
   FA_C_2_3_22 : FA_412 port map( A => q_2_3_22_port, B => q_2_4_22_port, Ci =>
                           q_2_5_22_port, S => q_3_2_22_port, Co => 
                           q_3_3_23_port, clk => clk);
   FA_C_2_3_23 : FA_411 port map( A => q_2_3_23_port, B => q_2_4_23_port, Ci =>
                           q_2_5_23_port, S => q_3_2_23_port, Co => 
                           q_3_3_24_port, clk => clk);
   FA_C_2_3_24 : FA_410 port map( A => q_2_3_24_port, B => q_2_4_24_port, Ci =>
                           q_2_5_24_port, S => q_3_2_24_port, Co => 
                           q_3_3_25_port, clk => clk);
   FA_C_2_3_25 : FA_409 port map( A => q_2_3_25_port, B => q_2_4_25_port, Ci =>
                           q_2_5_25_port, S => q_3_2_25_port, Co => 
                           q_3_3_26_port, clk => clk);
   FA_C_2_3_26 : FA_408 port map( A => q_2_3_26_port, B => q_2_4_26_port, Ci =>
                           q_2_5_26_port, S => q_3_2_26_port, Co => 
                           q_3_3_27_port, clk => clk);
   FA_C_2_3_27 : FA_407 port map( A => q_2_3_27_port, B => q_2_4_27_port, Ci =>
                           q_2_5_27_port, S => q_3_2_27_port, Co => 
                           q_3_3_28_port, clk => clk);
   FA_C_2_3_28 : FA_406 port map( A => q_2_3_28_port, B => q_2_4_28_port, Ci =>
                           q_2_5_28_port, S => q_3_2_28_port, Co => n366, clk 
                           => clk);
   FA_C_2_3_29 : FA_405 port map( A => q_2_3_29_port, B => q_2_4_29_port, Ci =>
                           q_2_5_29_port, S => q_3_2_29_port, Co => 
                           q_3_3_30_port, clk => clk);
   FA_C_2_3_30 : FA_404 port map( A => q_2_3_30_port, B => q_2_4_30_port, Ci =>
                           q_2_5_30_port, S => n369, Co => q_3_3_31_port, clk 
                           => clk);
   FA_C_2_3_31 : FA_403 port map( A => q_2_3_31_port, B => q_2_4_31_port, Ci =>
                           q_2_5_31_port, S => n371, Co => q_3_3_32_port, clk 
                           => clk);
   FA_C_2_3_32 : FA_402 port map( A => q_2_3_32_port, B => q_2_4_32_port, Ci =>
                           q_2_5_32_port, S => q_3_2_32_port, Co => 
                           q_3_3_33_port, clk => clk);
   FA_C_2_3_33 : FA_401 port map( A => n365, B => q_2_4_33_port, Ci => 
                           q_2_5_33_port, S => q_3_2_33_port, Co => 
                           q_3_3_34_port, clk => clk);
   FA_C_2_3_34 : FA_400 port map( A => q_2_3_34_port, B => q_2_4_34_port, Ci =>
                           q_2_5_34_port, S => q_3_2_34_port, Co => 
                           q_3_3_35_port, clk => clk);
   FA_C_2_3_35 : FA_399 port map( A => q_2_3_35_port, B => q_2_4_35_port, Ci =>
                           q_2_5_35_port, S => q_3_2_35_port, Co => 
                           q_3_3_36_port, clk => clk);
   FA_C_2_3_36 : FA_398 port map( A => q_2_3_36_port, B => q_2_4_36_port, Ci =>
                           q_2_5_36_port, S => q_3_2_36_port, Co => 
                           q_3_3_37_port, clk => clk);
   FA_C_2_3_37 : FA_397 port map( A => q_2_3_37_port, B => q_2_4_37_port, Ci =>
                           q_2_5_37_port, S => q_3_2_37_port, Co => 
                           q_3_3_38_port, clk => clk);
   FA_C_2_3_38 : FA_396 port map( A => q_2_3_38_port, B => q_2_4_38_port, Ci =>
                           q_2_5_38_port, S => q_3_2_38_port, Co => 
                           q_3_3_39_port, clk => clk);
   FA_C_2_3_39 : FA_395 port map( A => q_2_3_39_port, B => q_2_4_39_port, Ci =>
                           q_2_5_39_port, S => q_3_2_39_port, Co => 
                           q_3_3_40_port, clk => clk);
   FA_C_2_3_40 : FA_394 port map( A => q_2_3_40_port, B => q_2_4_40_port, Ci =>
                           q_2_5_40_port, S => q_3_2_40_port, Co => 
                           q_3_3_41_port, clk => clk);
   FA_C_2_3_41 : FA_393 port map( A => q_2_3_41_port, B => q_2_4_41_port, Ci =>
                           q_2_5_41_port, S => q_3_2_41_port, Co => 
                           q_3_3_42_port, clk => clk);
   FA_C_2_3_42 : FA_392 port map( A => q_2_3_42_port, B => q_2_4_42_port, Ci =>
                           q_2_5_42_port, S => q_3_2_42_port, Co => 
                           q_3_3_43_port, clk => clk);
   FA_C_2_3_43 : FA_391 port map( A => q_2_3_43_port, B => q_2_4_43_port, Ci =>
                           q_2_5_43_port, S => n364, Co => q_3_3_44_port, clk 
                           => clk);
   FA_C_2_3_44 : FA_390 port map( A => q_2_3_44_port, Ci => q_2_5_44_port, S =>
                           q_3_2_44_port, Co => q_3_3_45_port, B_BAR => 
                           q_2_4_44_port, clk => clk);
   FA_C_2_3_45 : FA_389 port map( A => q_2_3_45_port, Ci => q_2_5_45_port, S =>
                           q_3_2_45_port, Co => q_3_3_46_port, B_BAR => 
                           q_2_4_45_port, clk => clk);
   FA_C_2_3_46 : FA_388 port map( A => q_2_3_46_port, Ci => net102796, Co => 
                           q_3_3_47_port, B_BAR => q_2_4_46_port, S_BAR => 
                           q_3_2_46_port);
   FA_C_2_3_47 : FA_387 port map( A => q_2_3_47_port, B => net102794, Ci => 
                           net102795, S => q_3_2_47_port, Co => n_2039);
   HA_R_2_6_14 : HA_14 port map( A => q_0_6_14_port, B => q_0_7_14_port, S => 
                           q_3_4_14_port, C => q_3_5_15_port);
   HA_R_2_6_15 : HA_13 port map( A => q_0_6_15_port, B => q_0_7_15_port, S => 
                           q_3_4_15_port, C => q_3_5_16_port);
   FA_C_2_6_16 : FA_380 port map( A => q_0_7_16_port, B => q_0_8_16_port, Ci =>
                           B(17), S => q_3_4_16_port, Co => q_3_5_17_port);
   FA_C_2_6_17 : FA_379 port map( A => q_0_6_17_port, B => q_0_7_17_port, Ci =>
                           q_0_8_17_port, S => q_3_4_17_port, Co => 
                           q_3_5_18_port);
   FA_C_2_6_18 : FA_378 port map( A => q_0_8_18_port, B => q_0_9_18_port, S => 
                           q_3_4_18_port, Co => q_3_5_19_port, clk => clk, Ci 
                           => B(19));
   FA_C_2_6_19 : FA_377 port map( A => q_0_7_19_port, B => q_0_8_19_port, Ci =>
                           q_0_9_19_port, S => q_3_4_19_port, Co => 
                           q_3_5_20_port);
   FA_C_2_6_20 : FA_376 port map( A => q_0_9_20_port, B => q_0_10_20_port, Ci 
                           => B(21), S => q_3_4_20_port, Co => q_3_5_21_port);
   FA_C_2_6_21 : FA_375 port map( A => q_0_8_21_port, B => q_0_9_21_port, Ci =>
                           q_0_10_21_port, S => q_3_4_21_port, Co => 
                           q_3_5_22_port);
   FA_C_2_6_22 : FA_374 port map( A => q_2_6_22_port, B => q_0_11_22_port, Ci 
                           => n379, S => q_3_4_22_port, Co => q_3_5_23_port);
   FA_C_2_6_23 : FA_373 port map( A => n356, B => q_2_7_23_port, Ci => 
                           q_0_11_23_port, S => q_3_4_23_port, Co => 
                           q_3_5_24_port);
   FA_C_2_6_24 : FA_372 port map( A => q_2_6_24_port, B => q_2_7_24_port, Ci =>
                           n219, S => q_3_4_24_port, Co => q_3_5_25_port);
   FA_C_2_6_25 : FA_371 port map( A => q_2_6_25_port, B => q_2_7_25_port, Ci =>
                           q_0_12_25_port, S => q_3_4_25_port, Co => 
                           q_3_5_26_port, clk => clk);
   FA_C_2_6_26 : FA_370 port map( A => q_2_6_26_port, B => q_2_7_26_port, Ci =>
                           net102793, S => q_3_4_26_port, Co => q_3_5_27_port);
   FA_C_2_6_27 : FA_369 port map( A => q_2_6_27_port, B => q_2_7_27_port, Ci =>
                           net102792, S => q_3_4_27_port, Co => q_3_5_28_port);
   FA_C_2_6_28 : FA_368 port map( A => q_2_6_28_port, B => q_2_7_28_port, Ci =>
                           net102791, S => q_3_4_28_port, Co => q_3_5_29_port);
   FA_C_2_6_29 : FA_367 port map( A => q_2_6_29_port, B => net102789, Ci => 
                           net102790, S => q_3_4_29_port, Co => n_2040);
   FA_C_2_6_30 : FA_366 port map( A => net102787, B => q_2_7_30_port, Ci => 
                           net102788, S => q_3_4_30_port, Co => n_2041);
   FA_C_2_6_31 : FA_365 port map( B => net102785, Ci => net102786, Co => n_2042
                           , A_BAR => q_2_6_31_port, S_BAR => q_3_4_31_port);
   HA_R_3_0_6 : HA_11 port map( A => q_0_0_6_port, B => q_0_1_6_port, S => 
                           q_4_0_6_port, C => q_4_1_7_port);
   HA_R_3_0_7 : HA_10 port map( A => q_0_0_7_port, B => q_0_1_7_port, S => 
                           q_4_0_7_port, C => q_4_1_8_port);
   FA_C_3_0_8 : FA_344 port map( A => q_0_0_8_port, B => q_0_1_8_port, Ci => 
                           q_0_2_8_port, S => q_4_0_8_port, Co => q_4_1_9_port)
                           ;
   FA_C_3_0_9 : FA_343 port map( A => q_0_0_9_port, B => q_0_1_9_port, Ci => 
                           q_0_2_9_port, S => q_4_0_9_port, Co => q_4_1_10_port
                           );
   FA_C_3_0_10 : FA_342 port map( A => n355, B => q_0_2_10_port, Ci => 
                           q_0_3_10_port, S => q_4_0_10_port, Co => 
                           q_4_1_11_port);
   FA_C_3_0_11 : FA_341 port map( A => n354, B => q_3_1_11_port, Ci => 
                           q_0_2_11_port, S => q_4_0_11_port, Co => 
                           q_4_1_12_port);
   FA_C_3_0_12 : FA_340 port map( A => q_3_0_12_port, B => q_3_1_12_port, Ci =>
                           q_3_2_12_port, S => q_4_0_12_port, Co => 
                           q_4_1_13_port, clk => clk);
   FA_C_3_0_13 : FA_339 port map( A => q_3_0_13_port, B => q_3_1_13_port, Ci =>
                           q_3_2_13_port, S => q_4_0_13_port, Co => 
                           q_4_1_14_port, clk => clk);
   FA_C_3_0_14 : FA_338 port map( A => q_3_0_14_port, B => q_3_1_14_port, Ci =>
                           q_3_2_14_port, S => q_4_0_14_port, Co => 
                           q_4_1_15_port, clk => clk);
   FA_C_3_0_15 : FA_337 port map( A => q_3_0_15_port, B => q_3_1_15_port, Ci =>
                           q_3_2_15_port, S => q_4_0_15_port, Co => 
                           q_4_1_16_port, clk => clk);
   FA_C_3_0_16 : FA_336 port map( A => q_3_0_16_port, B => q_3_1_16_port, Ci =>
                           q_3_2_16_port, S => q_4_0_16_port, Co => 
                           q_4_1_17_port, clk => clk);
   FA_C_3_0_17 : FA_335 port map( A => q_3_0_17_port, B => q_3_1_17_port, Ci =>
                           q_3_2_17_port, S => q_4_0_17_port, Co => 
                           q_4_1_18_port, clk => clk);
   FA_C_3_0_18 : FA_334 port map( A => q_3_0_18_port, B => q_3_1_18_port, Ci =>
                           q_3_2_18_port, S => q_4_0_18_port, Co => 
                           q_4_1_19_port, clk => clk);
   FA_C_3_0_19 : FA_333 port map( A => q_3_0_19_port, B => q_3_1_19_port, Ci =>
                           q_3_2_19_port, S => q_4_0_19_port, Co => 
                           q_4_1_20_port, clk => clk);
   FA_C_3_0_20 : FA_332 port map( A => q_3_0_20_port, B => q_3_1_20_port, Ci =>
                           q_3_2_20_port, S => q_4_0_20_port, Co => 
                           q_4_1_21_port);
   FA_C_3_0_21 : FA_331 port map( A => q_3_0_21_port, B => q_3_1_21_port, Ci =>
                           n370, S => q_4_0_21_port, Co => q_4_1_22_port);
   FA_C_3_0_22 : FA_330 port map( A => q_3_0_22_port, B => q_3_1_22_port, Ci =>
                           q_3_2_22_port, S => q_4_0_22_port, Co => 
                           q_4_1_23_port);
   FA_C_3_0_23 : FA_329 port map( A => n373, B => q_3_1_23_port, Ci => 
                           q_3_2_23_port, S => q_4_0_23_port, Co => 
                           q_4_1_24_port, clk => clk);
   FA_C_3_0_24 : FA_328 port map( A => q_3_0_24_port, B => q_3_1_24_port, Ci =>
                           q_3_2_24_port, S => q_4_0_24_port, Co => 
                           q_4_1_25_port);
   FA_C_3_0_25 : FA_327 port map( A => q_3_0_25_port, B => q_3_1_25_port, Ci =>
                           q_3_2_25_port, S => q_4_0_25_port, Co => 
                           q_4_1_26_port);
   FA_C_3_0_26 : FA_326 port map( A => q_3_0_26_port, B => q_3_1_26_port, Ci =>
                           q_3_2_26_port, S => q_4_0_26_port, Co => n360);
   FA_C_3_0_27 : FA_325 port map( A => q_3_0_27_port, B => q_3_1_27_port, Ci =>
                           q_3_2_27_port, S => q_4_0_27_port, Co => 
                           q_4_1_28_port);
   FA_C_3_0_28 : FA_324 port map( A => q_3_0_28_port, B => q_3_1_28_port, Ci =>
                           q_3_2_28_port, S => q_4_0_28_port, Co => 
                           q_4_1_29_port);
   FA_C_3_0_29 : FA_323 port map( A => q_3_0_29_port, B => q_3_1_29_port, Ci =>
                           q_3_2_29_port, S => n359, Co => q_4_1_30_port);
   FA_C_3_0_30 : FA_322 port map( A => q_3_0_30_port, B => q_3_1_30_port, Ci =>
                           n369, S => q_4_0_30_port, Co => q_4_1_31_port);
   FA_C_3_0_31 : FA_321 port map( A => q_3_0_31_port, B => q_3_1_31_port, Ci =>
                           n371, S => q_4_0_31_port, Co => q_4_1_32_port);
   FA_C_3_0_32 : FA_320 port map( A => q_3_0_32_port, B => q_3_1_32_port, Ci =>
                           q_3_2_32_port, S => q_4_0_32_port, Co => 
                           q_4_1_33_port);
   FA_C_3_0_33 : FA_319 port map( A => q_3_0_33_port, B => q_3_1_33_port, Ci =>
                           q_3_2_33_port, S => q_4_0_33_port, Co => 
                           q_4_1_34_port);
   FA_C_3_0_34 : FA_318 port map( A => q_3_0_34_port, B => q_3_1_34_port, Ci =>
                           q_3_2_34_port, S => n349, Co => q_4_1_35_port);
   FA_C_3_0_35 : FA_317 port map( A => q_3_0_35_port, B => n353, Ci => 
                           q_3_2_35_port, S => n346, Co => q_4_1_36_port);
   FA_C_3_0_36 : FA_316 port map( A => q_3_0_36_port, B => q_3_1_36_port, Ci =>
                           q_3_2_36_port, S => q_4_0_36_port, Co => 
                           q_4_1_37_port);
   FA_C_3_0_37 : FA_315 port map( A => q_3_0_37_port, B => q_3_1_37_port, Ci =>
                           q_3_2_37_port, S => q_4_0_37_port, Co => 
                           q_4_1_38_port);
   FA_C_3_0_38 : FA_314 port map( A => q_3_0_38_port, B => q_3_1_38_port, Ci =>
                           q_3_2_38_port, S => q_4_0_38_port, Co => 
                           q_4_1_39_port);
   FA_C_3_0_39 : FA_313 port map( A => q_3_0_39_port, B => q_3_1_39_port, Ci =>
                           q_3_2_39_port, S => q_4_0_39_port, Co => 
                           q_4_1_40_port);
   FA_C_3_0_40 : FA_312 port map( A => q_3_0_40_port, B => q_3_1_40_port, Ci =>
                           q_3_2_40_port, S => q_4_0_40_port, Co => 
                           q_4_1_41_port);
   FA_C_3_0_41 : FA_311 port map( A => q_3_0_41_port, B => q_3_1_41_port, Ci =>
                           q_3_2_41_port, S => q_4_0_41_port, Co => 
                           q_4_1_42_port);
   FA_C_3_0_42 : FA_310 port map( A => q_3_0_42_port, B => q_3_1_42_port, Ci =>
                           q_3_2_42_port, S => q_4_0_42_port, Co => 
                           q_4_1_43_port);
   FA_C_3_0_43 : FA_309 port map( A => n367, B => q_3_1_43_port, Ci => n364, S 
                           => q_4_0_43_port, Co => q_4_1_44_port);
   FA_C_3_0_44 : FA_308 port map( A => q_3_0_44_port, B => n368, Ci => 
                           q_3_2_44_port, S => q_4_0_44_port, Co => 
                           q_4_1_45_port);
   FA_C_3_0_45 : FA_307 port map( A => q_3_0_45_port, B => q_3_1_45_port, Ci =>
                           q_3_2_45_port, S => q_4_0_45_port, Co => 
                           q_4_1_46_port);
   FA_C_3_0_46 : FA_306 port map( A => q_3_0_46_port, B => q_3_1_46_port, S => 
                           q_4_0_46_port, Co => q_4_1_47_port, Ci_BAR => 
                           q_3_2_46_port, clk => clk);
   FA_C_3_0_47 : FA_305 port map( A => q_3_0_47_port, B => q_3_1_47_port, Ci =>
                           q_3_2_47_port, S => q_4_0_47_port, Co => n_2043, clk
                           => clk);
   HA_R_3_3_8 : HA_8 port map( A => q_0_3_8_port, B => q_0_4_8_port, S => 
                           q_4_2_8_port, C => q_5_2_9_port);
   HA_R_3_3_9 : HA_7 port map( A => q_0_3_9_port, B => q_0_4_9_port, S => 
                           q_4_2_9_port, C => q_5_2_10_port);
   FA_C_3_3_10 : FA_292 port map( A => q_0_4_10_port, B => q_0_5_10_port, S => 
                           q_4_2_10_port, Co => q_5_2_11_port, Ci_BAR => n230);
   FA_C_3_3_11 : FA_291 port map( A => q_0_3_11_port, B => q_0_4_11_port, Ci =>
                           q_0_5_11_port, S => q_4_2_11_port, Co => 
                           q_5_2_12_port);
   FA_C_3_3_12 : FA_290 port map( A => q_0_5_12_port, B => q_0_6_12_port, Ci =>
                           B(13), S => q_4_2_12_port, Co => q_5_2_13_port);
   FA_C_3_3_13 : FA_289 port map( A => q_3_3_13_port, B => q_0_5_13_port, Ci =>
                           q_0_6_13_port, S => q_4_2_13_port, Co => 
                           q_5_2_14_port, clk => clk);
   FA_C_3_3_14 : FA_288 port map( A => q_3_3_14_port, B => q_3_4_14_port, S => 
                           q_4_2_14_port, Co => q_5_2_15_port, Ci => B(15), clk
                           => clk);
   FA_C_3_3_15 : FA_287 port map( A => q_3_3_15_port, B => q_3_4_15_port, Ci =>
                           q_3_5_15_port, S => q_4_2_15_port, Co => 
                           q_5_2_16_port, clk => clk);
   FA_C_3_3_16 : FA_286 port map( A => q_3_3_16_port, B => q_3_4_16_port, Ci =>
                           q_3_5_16_port, S => q_4_2_16_port, Co => 
                           q_5_2_17_port, clk => clk);
   FA_C_3_3_17 : FA_285 port map( A => q_3_3_17_port, B => q_3_4_17_port, Ci =>
                           q_3_5_17_port, S => q_4_2_17_port, Co => 
                           q_5_2_18_port, clk => clk);
   FA_C_3_3_18 : FA_284 port map( A => q_3_3_18_port, B => q_3_4_18_port, Ci =>
                           q_3_5_18_port, S => q_4_2_18_port, Co => 
                           q_5_2_19_port, clk => clk);
   FA_C_3_3_19 : FA_283 port map( A => q_3_3_19_port, B => q_3_4_19_port, Ci =>
                           q_3_5_19_port, S => q_4_2_19_port, Co => 
                           q_5_2_20_port, clk => clk);
   FA_C_3_3_20 : FA_282 port map( A => q_3_3_20_port, B => q_3_4_20_port, Ci =>
                           q_3_5_20_port, S => q_4_2_20_port, Co => 
                           q_5_2_21_port, clk => clk);
   FA_C_3_3_21 : FA_281 port map( A => q_3_3_21_port, B => q_3_4_21_port, Ci =>
                           q_3_5_21_port, S => q_4_2_21_port, Co => 
                           q_5_2_22_port, clk => clk);
   FA_C_3_3_22 : FA_280 port map( A => q_3_3_22_port, B => q_3_4_22_port, Ci =>
                           q_3_5_22_port, S => q_4_2_22_port, Co => 
                           q_5_2_23_port, clk => clk);
   FA_C_3_3_23 : FA_279 port map( A => q_3_3_23_port, B => q_3_4_23_port, Ci =>
                           q_3_5_23_port, S => q_4_2_23_port, Co => 
                           q_5_2_24_port, clk => clk);
   FA_C_3_3_24 : FA_278 port map( A => q_3_3_24_port, B => q_3_4_24_port, Ci =>
                           q_3_5_24_port, S => q_4_2_24_port, Co => 
                           q_5_2_25_port, clk => clk);
   FA_C_3_3_25 : FA_277 port map( A => q_3_3_25_port, B => q_3_4_25_port, Ci =>
                           q_3_5_25_port, S => q_4_2_25_port, Co => 
                           q_5_2_26_port, clk => clk);
   FA_C_3_3_26 : FA_276 port map( A => q_3_3_26_port, B => q_3_4_26_port, Ci =>
                           q_3_5_26_port, S => q_4_2_26_port, Co => 
                           q_5_2_27_port, clk => clk);
   FA_C_3_3_27 : FA_275 port map( A => q_3_3_27_port, B => q_3_4_27_port, Ci =>
                           q_3_5_27_port, S => q_4_2_27_port, Co => 
                           q_5_2_28_port, clk => clk);
   FA_C_3_3_28 : FA_274 port map( A => q_3_3_28_port, B => q_3_4_28_port, Ci =>
                           q_3_5_28_port, S => q_4_2_28_port, Co => 
                           q_5_2_29_port, clk => clk);
   FA_C_3_3_29 : FA_273 port map( A => n366, B => q_3_4_29_port, Ci => 
                           q_3_5_29_port, S => n358, Co => q_5_2_30_port, clk 
                           => clk);
   FA_C_3_3_30 : FA_272 port map( A => q_3_3_30_port, B => q_3_4_30_port, Ci =>
                           net102784, S => q_4_2_30_port, Co => q_5_2_31_port, 
                           clk => clk);
   FA_C_3_3_31 : FA_271 port map( A => q_3_3_31_port, Ci => net102783, S => 
                           q_4_2_31_port, Co => q_5_2_32_port, B_BAR => 
                           q_3_4_31_port, clk => clk);
   FA_C_3_3_32 : FA_270 port map( A => q_3_3_32_port, B => net102781, Ci => 
                           net102782, S => q_4_2_32_port, Co => n_2044);
   FA_C_3_3_33 : FA_269 port map( A => q_3_3_33_port, B => net102779, Ci => 
                           net102780, S => q_4_2_33_port, Co => n_2045);
   FA_C_3_3_34 : FA_268 port map( A => q_3_3_34_port, B => net102777, Ci => 
                           net102778, S => q_4_2_34_port, Co => n_2046);
   FA_C_3_3_35 : FA_267 port map( A => q_3_3_35_port, B => net102775, Ci => 
                           net102776, S => q_4_2_35_port, Co => n_2047);
   FA_C_3_3_36 : FA_266 port map( A => q_3_3_36_port, B => net102773, Ci => 
                           net102774, S => q_4_2_36_port, Co => n_2048);
   FA_C_3_3_37 : FA_265 port map( A => q_3_3_37_port, B => net102771, Ci => 
                           net102772, S => q_4_2_37_port, Co => n_2049);
   FA_C_3_3_38 : FA_264 port map( A => q_3_3_38_port, B => net102769, Ci => 
                           net102770, S => q_4_2_38_port, Co => n_2050);
   FA_C_3_3_39 : FA_263 port map( A => q_3_3_39_port, B => net102767, Ci => 
                           net102768, S => q_4_2_39_port, Co => n_2051);
   FA_C_3_3_40 : FA_262 port map( A => q_3_3_40_port, B => net102765, Ci => 
                           net102766, S => q_4_2_40_port, Co => n_2052);
   FA_C_3_3_41 : FA_261 port map( A => q_3_3_41_port, B => net102763, Ci => 
                           net102764, S => q_4_2_41_port, Co => n_2053);
   FA_C_3_3_42 : FA_260 port map( A => q_3_3_42_port, B => net102761, Ci => 
                           net102762, S => q_4_2_42_port, Co => n_2054);
   FA_C_3_3_43 : FA_259 port map( A => q_3_3_43_port, B => net102759, Ci => 
                           net102760, S => q_4_2_43_port, Co => n_2055);
   FA_C_3_3_44 : FA_258 port map( A => q_3_3_44_port, B => net102757, Ci => 
                           net102758, S => q_4_2_44_port, Co => n_2056);
   FA_C_3_3_45 : FA_257 port map( A => q_3_3_45_port, B => net102755, Ci => 
                           net102756, S => q_4_2_45_port, Co => n_2057);
   FA_C_3_3_46 : FA_256 port map( A => q_3_3_46_port, B => net102753, Ci => 
                           net102754, S => q_4_2_46_port, Co => n_2058);
   FA_C_3_3_47 : FA_255 port map( A => q_3_3_47_port, B => net102751, Ci => 
                           net102752, S => q_4_2_47_port, Co => n_2059);
   HA_R_4_0_4 : HA_5 port map( A => q_0_0_4_port, B => q_0_1_4_port, S => 
                           q_5_0_4_port, C => q_5_1_5_port);
   HA_R_4_0_5 : HA_4 port map( A => q_0_0_5_port, B => q_0_1_5_port, S => 
                           q_5_0_5_port, C => q_5_1_6_port);
   FA_C_4_0_6 : FA_244 port map( A => q_4_0_6_port, B => q_0_2_6_port, Ci => 
                           q_0_3_6_port, S => q_5_0_6_port, Co => n376, clk => 
                           clk);
   FA_C_4_0_7 : FA_243 port map( A => q_4_0_7_port, B => q_4_1_7_port, Ci => 
                           q_0_2_7_port, S => n375, Co => q_5_1_8_port, clk => 
                           clk);
   FA_C_4_0_8 : FA_242 port map( A => q_4_0_8_port, B => q_4_1_8_port, Ci => 
                           q_4_2_8_port, S => q_5_0_8_port, Co => q_5_1_9_port,
                           clk => clk);
   FA_C_4_0_9 : FA_241 port map( A => q_4_0_9_port, B => q_4_1_9_port, Ci => 
                           q_4_2_9_port, S => q_5_0_9_port, Co => q_5_1_10_port
                           , clk => clk);
   FA_C_4_0_10 : FA_240 port map( A => q_4_0_10_port, B => q_4_1_10_port, Ci =>
                           q_4_2_10_port, S => q_5_0_10_port, Co => 
                           q_5_1_11_port, clk => clk);
   FA_C_4_0_11 : FA_239 port map( A => q_4_0_11_port, B => q_4_1_11_port, Ci =>
                           q_4_2_11_port, S => q_5_0_11_port, Co => 
                           q_5_1_12_port, clk => clk);
   FA_C_4_0_12 : FA_238 port map( A => q_4_0_12_port, B => q_4_1_12_port, Ci =>
                           q_4_2_12_port, S => q_5_0_12_port, Co => 
                           q_5_1_13_port, clk => clk);
   FA_C_4_0_13 : FA_237 port map( A => q_4_0_13_port, B => q_4_1_13_port, Ci =>
                           q_4_2_13_port, S => q_5_0_13_port, Co => 
                           q_5_1_14_port);
   FA_C_4_0_14 : FA_236 port map( A => q_4_0_14_port, B => q_4_1_14_port, Ci =>
                           q_4_2_14_port, S => q_5_0_14_port, Co => 
                           q_5_1_15_port, clk => clk);
   FA_C_4_0_15 : FA_235 port map( A => q_4_0_15_port, B => q_4_1_15_port, Ci =>
                           q_4_2_15_port, S => q_5_0_15_port, Co => 
                           q_5_1_16_port);
   FA_C_4_0_16 : FA_234 port map( A => q_4_0_16_port, B => q_4_1_16_port, Ci =>
                           q_4_2_16_port, S => q_5_0_16_port, Co => 
                           q_5_1_17_port);
   FA_C_4_0_17 : FA_233 port map( A => q_4_0_17_port, B => q_4_1_17_port, Ci =>
                           q_4_2_17_port, S => q_5_0_17_port, Co => 
                           q_5_1_18_port);
   FA_C_4_0_18 : FA_232 port map( A => q_4_0_18_port, B => q_4_1_18_port, Ci =>
                           q_4_2_18_port, S => q_5_0_18_port, Co => 
                           q_5_1_19_port);
   FA_C_4_0_19 : FA_231 port map( A => q_4_0_19_port, B => q_4_1_19_port, Ci =>
                           q_4_2_19_port, S => q_5_0_19_port, Co => 
                           q_5_1_20_port);
   FA_C_4_0_20 : FA_230 port map( A => q_4_0_20_port, B => q_4_1_20_port, Ci =>
                           q_4_2_20_port, S => q_5_0_20_port, Co => 
                           q_5_1_21_port);
   FA_C_4_0_21 : FA_229 port map( A => q_4_0_21_port, B => q_4_1_21_port, Ci =>
                           q_4_2_21_port, S => q_5_0_21_port, Co => n343);
   FA_C_4_0_22 : FA_228 port map( A => q_4_0_22_port, B => q_4_1_22_port, Ci =>
                           q_4_2_22_port, S => q_5_0_22_port, Co => 
                           q_5_1_23_port);
   FA_C_4_0_23 : FA_227 port map( A => q_4_0_23_port, B => q_4_1_23_port, Ci =>
                           q_4_2_23_port, S => q_5_0_23_port, Co => 
                           q_5_1_24_port);
   FA_C_4_0_24 : FA_226 port map( A => q_4_0_24_port, B => q_4_1_24_port, Ci =>
                           q_4_2_24_port, S => q_5_0_24_port, Co => 
                           q_5_1_25_port);
   FA_C_4_0_25 : FA_225 port map( A => q_4_0_25_port, B => q_4_1_25_port, Ci =>
                           q_4_2_25_port, S => q_5_0_25_port, Co => 
                           q_5_1_26_port);
   FA_C_4_0_26 : FA_224 port map( A => q_4_0_26_port, B => q_4_1_26_port, Ci =>
                           q_4_2_26_port, S => q_5_0_26_port, Co => 
                           q_5_1_27_port);
   FA_C_4_0_27 : FA_223 port map( A => q_4_0_27_port, B => n360, Ci => 
                           q_4_2_27_port, S => n345, Co => n344);
   FA_C_4_0_28 : FA_222 port map( A => q_4_0_28_port, B => q_4_1_28_port, Ci =>
                           q_4_2_28_port, S => q_5_0_28_port, Co => 
                           q_5_1_29_port);
   FA_C_4_0_29 : FA_221 port map( A => n359, B => q_4_1_29_port, Ci => n358, S 
                           => q_5_0_29_port, Co => q_5_1_30_port);
   FA_C_4_0_30 : FA_220 port map( A => q_4_0_30_port, B => q_4_1_30_port, Ci =>
                           q_4_2_30_port, S => q_5_0_30_port, Co => 
                           q_5_1_31_port);
   FA_C_4_0_31 : FA_219 port map( A => q_4_0_31_port, B => q_4_1_31_port, Ci =>
                           q_4_2_31_port, S => q_5_0_31_port, Co => 
                           q_5_1_32_port);
   FA_C_4_0_32 : FA_218 port map( A => q_4_0_32_port, B => q_4_1_32_port, S => 
                           q_5_0_32_port, Co => q_5_1_33_port, Ci => 
                           q_4_2_32_port);
   FA_C_4_0_33 : FA_217 port map( A => q_4_0_33_port, B => q_4_1_33_port, Ci =>
                           q_4_2_33_port, S => q_5_0_33_port, Co => 
                           q_5_1_34_port);
   FA_C_4_0_34 : FA_216 port map( A => n349, B => q_4_1_34_port, S => 
                           q_5_0_34_port, Co => q_5_1_35_port, Ci => 
                           q_4_2_34_port);
   FA_C_4_0_35 : FA_215 port map( A => n346, B => q_4_1_35_port, Ci => 
                           q_4_2_35_port, S => q_5_0_35_port, Co => 
                           q_5_1_36_port);
   FA_C_4_0_36 : FA_214 port map( A => q_4_0_36_port, B => q_4_1_36_port, Ci =>
                           q_4_2_36_port, S => q_5_0_36_port, Co => 
                           q_5_1_37_port);
   FA_C_4_0_37 : FA_213 port map( A => q_4_0_37_port, B => q_4_1_37_port, Ci =>
                           q_4_2_37_port, S => q_5_0_37_port, Co => 
                           q_5_1_38_port);
   FA_C_4_0_38 : FA_212 port map( A => q_4_0_38_port, B => q_4_1_38_port, Ci =>
                           q_4_2_38_port, S => q_5_0_38_port, Co => 
                           q_5_1_39_port);
   FA_C_4_0_39 : FA_211 port map( A => q_4_0_39_port, B => q_4_1_39_port, S => 
                           q_5_0_39_port, Co => q_5_1_40_port, Ci => 
                           q_4_2_39_port);
   FA_C_4_0_40 : FA_210 port map( A => q_4_0_40_port, B => q_4_1_40_port, Ci =>
                           q_4_2_40_port, S => q_5_0_40_port, Co => 
                           q_5_1_41_port);
   FA_C_4_0_41 : FA_209 port map( A => q_4_0_41_port, B => q_4_1_41_port, Ci =>
                           q_4_2_41_port, S => q_5_0_41_port, Co => 
                           q_5_1_42_port);
   FA_C_4_0_42 : FA_208 port map( A => q_4_0_42_port, B => q_4_1_42_port, Ci =>
                           q_4_2_42_port, S => q_5_0_42_port, Co => 
                           q_5_1_43_port);
   FA_C_4_0_43 : FA_207 port map( A => q_4_0_43_port, B => q_4_1_43_port, Ci =>
                           q_4_2_43_port, S => q_5_0_43_port, Co => n350);
   FA_C_4_0_44 : FA_206 port map( A => q_4_0_44_port, B => q_4_1_44_port, Ci =>
                           q_4_2_44_port, S => q_5_0_44_port, Co => 
                           q_5_1_45_port);
   FA_C_4_0_45 : FA_205 port map( A => q_4_0_45_port, B => q_4_1_45_port, S => 
                           q_5_0_45_port, Co => q_5_1_46_port, Ci => 
                           q_4_2_45_port);
   FA_C_4_0_46 : FA_204 port map( A => q_4_0_46_port, B => q_4_1_46_port, S => 
                           q_5_0_46_port, Co => q_5_1_47_port, Ci => 
                           q_4_2_46_port);
   FA_C_4_0_47 : FA_203 port map( A => q_4_0_47_port, B => q_4_1_47_port, Ci =>
                           q_4_2_47_port, S => q_5_0_47_port, Co => n_2060, clk
                           => clk);
   HA_R_5_0_2 : HA_2 port map( A => q_0_0_2_port, B => q_0_1_2_port, S => 
                           q_6_0_2_port, C => q_6_1_3_port);
   HA_R_5_0_3 : HA_1 port map( A => q_0_0_3_port, B => q_0_1_3_port, S => 
                           q_6_0_3_port, C => q_6_1_4_port);
   FA_C_5_0_4 : FA_188 port map( A => q_5_0_4_port, B => q_0_2_4_port, Ci => 
                           B(5), S => q_6_0_4_port, Co => q_6_1_5_port, clk => 
                           clk);
   FA_C_5_0_5 : FA_187 port map( A => q_5_0_5_port, B => q_5_1_5_port, Ci => 
                           q_0_2_5_port, S => q_6_0_5_port, Co => q_6_1_6_port,
                           clk => clk);
   FA_C_5_0_6 : FA_186 port map( A => q_5_0_6_port, B => q_5_1_6_port, S => 
                           q_6_0_6_port, Co => q_6_1_7_port, Ci_BAR => n227, 
                           clk => clk);
   FA_C_5_0_7 : FA_185 port map( A => n375, B => n376, Ci => q_0_3_7_port, S =>
                           q_6_0_7_port, Co => q_6_1_8_port, clk => clk);
   FA_C_5_0_8 : FA_184 port map( A => q_5_0_8_port, B => q_5_1_8_port, Ci => 
                           B(9), S => q_6_0_8_port, Co => q_6_1_9_port, clk => 
                           clk);
   FA_C_5_0_9 : FA_183 port map( A => q_5_0_9_port, B => q_5_1_9_port, Ci => 
                           q_5_2_9_port, S => q_6_0_9_port, Co => q_6_1_10_port
                           , clk => clk);
   FA_C_5_0_10 : FA_182 port map( A => q_5_0_10_port, B => q_5_1_10_port, Ci =>
                           q_5_2_10_port, S => q_6_0_10_port, Co => 
                           q_6_1_11_port, clk => clk);
   FA_C_5_0_11 : FA_181 port map( A => q_5_0_11_port, B => q_5_1_11_port, Ci =>
                           q_5_2_11_port, S => q_6_0_11_port, Co => 
                           q_6_1_12_port, clk => clk);
   FA_C_5_0_12 : FA_180 port map( A => q_5_0_12_port, B => q_5_1_12_port, Ci =>
                           q_5_2_12_port, S => q_6_0_12_port, Co => 
                           q_6_1_13_port, clk => clk);
   FA_C_5_0_13 : FA_179 port map( A => q_5_0_13_port, B => q_5_1_13_port, Ci =>
                           q_5_2_13_port, S => q_6_0_13_port, Co => 
                           q_6_1_14_port, clk => clk);
   FA_C_5_0_14 : FA_178 port map( A => q_5_0_14_port, B => q_5_1_14_port, Ci =>
                           q_5_2_14_port, S => q_6_0_14_port, Co => 
                           q_6_1_15_port, clk => clk);
   FA_C_5_0_15 : FA_177 port map( A => q_5_0_15_port, B => q_5_1_15_port, Ci =>
                           q_5_2_15_port, S => q_6_0_15_port, Co => 
                           q_6_1_16_port);
   FA_C_5_0_16 : FA_176 port map( A => q_5_0_16_port, B => q_5_1_16_port, Ci =>
                           q_5_2_16_port, S => q_6_0_16_port, Co => 
                           q_6_1_17_port);
   FA_C_5_0_17 : FA_175 port map( A => q_5_0_17_port, B => q_5_1_17_port, Ci =>
                           q_5_2_17_port, S => q_6_0_17_port, Co => 
                           q_6_1_18_port);
   FA_C_5_0_18 : FA_174 port map( A => q_5_0_18_port, B => q_5_1_18_port, Ci =>
                           q_5_2_18_port, S => q_6_0_18_port, Co => 
                           q_6_1_19_port);
   FA_C_5_0_19 : FA_173 port map( A => q_5_0_19_port, B => q_5_1_19_port, Ci =>
                           q_5_2_19_port, S => q_6_0_19_port, Co => 
                           q_6_1_20_port);
   FA_C_5_0_20 : FA_172 port map( A => q_5_0_20_port, B => q_5_1_20_port, Ci =>
                           q_5_2_20_port, S => q_6_0_20_port, Co => 
                           q_6_1_21_port);
   FA_C_5_0_21 : FA_171 port map( A => q_5_0_21_port, B => q_5_1_21_port, Ci =>
                           q_5_2_21_port, S => q_6_0_21_port, Co => 
                           q_6_1_22_port);
   FA_C_5_0_22 : FA_170 port map( A => q_5_0_22_port, B => n343, Ci => 
                           q_5_2_22_port, S => q_6_0_22_port, Co => 
                           q_6_1_23_port);
   FA_C_5_0_23 : FA_169 port map( A => q_5_0_23_port, B => q_5_1_23_port, Ci =>
                           q_5_2_23_port, S => q_6_0_23_port, Co => 
                           q_6_1_24_port);
   FA_C_5_0_24 : FA_168 port map( A => q_5_0_24_port, B => q_5_1_24_port, Ci =>
                           q_5_2_24_port, S => q_6_0_24_port, Co => 
                           q_6_1_25_port);
   FA_C_5_0_25 : FA_167 port map( A => q_5_0_25_port, B => q_5_1_25_port, Ci =>
                           q_5_2_25_port, S => q_6_0_25_port, Co => 
                           q_6_1_26_port);
   FA_C_5_0_26 : FA_166 port map( A => q_5_0_26_port, B => q_5_1_26_port, Ci =>
                           q_5_2_26_port, S => q_6_0_26_port, Co => 
                           q_6_1_27_port);
   FA_C_5_0_27 : FA_165 port map( A => n345, B => q_5_1_27_port, Ci => 
                           q_5_2_27_port, S => q_6_0_27_port, Co => 
                           q_6_1_28_port);
   FA_C_5_0_28 : FA_164 port map( A => q_5_0_28_port, B => n344, Ci => 
                           q_5_2_28_port, S => q_6_0_28_port, Co => 
                           q_6_1_29_port);
   FA_C_5_0_29 : FA_163 port map( A => q_5_0_29_port, B => q_5_1_29_port, Ci =>
                           q_5_2_29_port, S => q_6_0_29_port, Co => 
                           q_6_1_30_port);
   FA_C_5_0_30 : FA_162 port map( A => q_5_0_30_port, B => q_5_1_30_port, Ci =>
                           q_5_2_30_port, S => q_6_0_30_port, Co => 
                           q_6_1_31_port);
   FA_C_5_0_31 : FA_161 port map( A => q_5_0_31_port, B => q_5_1_31_port, Ci =>
                           q_5_2_31_port, S => q_6_0_31_port, Co => 
                           q_6_1_32_port, clk => clk);
   FA_C_5_0_32 : FA_160 port map( A => q_5_0_32_port, B => q_5_1_32_port, Ci =>
                           q_5_2_32_port, S => q_6_0_32_port, Co => 
                           q_6_1_33_port, clk => clk);
   FA_C_5_0_33 : FA_159 port map( A => q_5_0_33_port, B => q_5_1_33_port, Ci =>
                           net102750, S => q_6_0_33_port, Co => q_6_1_34_port);
   FA_C_5_0_34 : FA_158 port map( A => q_5_0_34_port, B => q_5_1_34_port, Ci =>
                           net102749, S => q_6_0_34_port, Co => q_6_1_35_port, 
                           clk => clk);
   FA_C_5_0_35 : FA_157 port map( A => q_5_0_35_port, B => q_5_1_35_port, Ci =>
                           net102748, S => q_6_0_35_port, Co => q_6_1_36_port, 
                           clk => clk);
   FA_C_5_0_36 : FA_156 port map( A => q_5_0_36_port, B => q_5_1_36_port, Ci =>
                           net102747, S => q_6_0_36_port, Co => n342, clk => 
                           clk);
   FA_C_5_0_37 : FA_155 port map( A => q_5_0_37_port, B => q_5_1_37_port, Ci =>
                           net102746, S => q_6_0_37_port, Co => q_6_1_38_port, 
                           clk => clk);
   FA_C_5_0_38 : FA_154 port map( A => q_5_0_38_port, B => q_5_1_38_port, Ci =>
                           net102745, S => q_6_0_38_port, Co => q_6_1_39_port, 
                           clk => clk);
   FA_C_5_0_39 : FA_153 port map( A => q_5_0_39_port, B => q_5_1_39_port, Ci =>
                           net102744, S => q_6_0_39_port, Co => q_6_1_40_port, 
                           clk => clk);
   FA_C_5_0_40 : FA_152 port map( A => q_5_0_40_port, B => q_5_1_40_port, Ci =>
                           net102743, S => q_6_0_40_port, Co => q_6_1_41_port, 
                           clk => clk);
   FA_C_5_0_41 : FA_151 port map( A => q_5_0_41_port, B => q_5_1_41_port, Ci =>
                           net102742, S => q_6_0_41_port, Co => q_6_1_42_port, 
                           clk => clk);
   FA_C_5_0_42 : FA_150 port map( A => q_5_0_42_port, B => q_5_1_42_port, Ci =>
                           net102741, S => q_6_0_42_port, Co => q_6_1_43_port, 
                           clk => clk);
   FA_C_5_0_43 : FA_149 port map( A => q_5_0_43_port, B => q_5_1_43_port, Ci =>
                           net102740, S => q_6_0_43_port, Co => q_6_1_44_port);
   FA_C_5_0_44 : FA_148 port map( A => q_5_0_44_port, B => n350, Ci => 
                           net102739, S => q_6_0_44_port, Co => q_6_1_45_port);
   FA_C_5_0_45 : FA_147 port map( A => q_5_0_45_port, B => q_5_1_45_port, Ci =>
                           net102738, S => q_6_0_45_port, Co => q_6_1_46_port);
   FA_C_5_0_46 : FA_146 port map( A => q_5_0_46_port, B => q_5_1_46_port, Ci =>
                           net102737, S => q_6_0_46_port, Co => q_6_1_47_port);
   FA_C_5_0_47 : FA_145 port map( A => q_5_0_47_port, B => q_5_1_47_port, Ci =>
                           net102736, S => q_6_0_47_port, Co => n_2061);
   P4_ADDER_0 : P4_ADDER_NBIT64_NBIT_PER_BLOCK4_NBLOCKS16 port map( A(63) => 
                           n182, A(62) => n183, A(61) => n184, A(60) => n185, 
                           A(59) => n186, A(58) => n187, A(57) => n188, A(56) 
                           => n189, A(55) => n190, A(54) => n191, A(53) => n192
                           , A(52) => n193, A(51) => n194, A(50) => n195, A(49)
                           => n196, A(48) => n197, A(47) => q_6_0_47_port, 
                           A(46) => q_6_0_46_port, A(45) => q_6_0_45_port, 
                           A(44) => q_6_0_44_port, A(43) => q_6_0_43_port, 
                           A(42) => q_6_0_42_port, A(41) => q_6_0_41_port, 
                           A(40) => q_6_0_40_port, A(39) => q_6_0_39_port, 
                           A(38) => q_6_0_38_port, A(37) => q_6_0_37_port, 
                           A(36) => q_6_0_36_port, A(35) => q_6_0_35_port, 
                           A(34) => q_6_0_34_port, A(33) => q_6_0_33_port, 
                           A(32) => q_6_0_32_port, A(31) => q_6_0_31_port, 
                           A(30) => q_6_0_30_port, A(29) => q_6_0_29_port, 
                           A(28) => q_6_0_28_port, A(27) => q_6_0_27_port, 
                           A(26) => q_6_0_26_port, A(25) => q_6_0_25_port, 
                           A(24) => q_6_0_24_port, A(23) => q_6_0_23_port, 
                           A(22) => q_6_0_22_port, A(21) => q_6_0_21_port, 
                           A(20) => q_6_0_20_port, A(19) => q_6_0_19_port, 
                           A(18) => q_6_0_18_port, A(17) => q_6_0_17_port, 
                           A(16) => q_6_0_16_port, A(15) => q_6_0_15_port, 
                           A(14) => q_6_0_14_port, A(13) => q_6_0_13_port, 
                           A(12) => q_6_0_12_port, A(11) => q_6_0_11_port, 
                           A(10) => q_6_0_10_port, A(9) => q_6_0_9_port, A(8) 
                           => q_6_0_8_port, A(7) => q_6_0_7_port, A(6) => 
                           q_6_0_6_port, A(5) => q_6_0_5_port, A(4) => 
                           q_6_0_4_port, A(3) => q_6_0_3_port, A(2) => 
                           q_6_0_2_port, A(1) => q_0_0_1_port, A(0) => 
                           q_0_0_0_port, B(63) => n198, B(62) => n199, B(61) =>
                           n200, B(60) => n201, B(59) => n202, B(58) => n203, 
                           B(57) => n204, B(56) => n205, B(55) => n206, B(54) 
                           => n207, B(53) => n208, B(52) => n209, B(51) => n210
                           , B(50) => n211, B(49) => n212, B(48) => n213, B(47)
                           => q_6_1_47_port, B(46) => q_6_1_46_port, B(45) => 
                           q_6_1_45_port, B(44) => q_6_1_44_port, B(43) => 
                           q_6_1_43_port, B(42) => q_6_1_42_port, B(41) => 
                           q_6_1_41_port, B(40) => q_6_1_40_port, B(39) => 
                           q_6_1_39_port, B(38) => q_6_1_38_port, B(37) => n342
                           , B(36) => q_6_1_36_port, B(35) => q_6_1_35_port, 
                           B(34) => q_6_1_34_port, B(33) => q_6_1_33_port, 
                           B(32) => q_6_1_32_port, B(31) => q_6_1_31_port, 
                           B(30) => q_6_1_30_port, B(29) => q_6_1_29_port, 
                           B(28) => q_6_1_28_port, B(27) => q_6_1_27_port, 
                           B(26) => q_6_1_26_port, B(25) => q_6_1_25_port, 
                           B(24) => q_6_1_24_port, B(23) => q_6_1_23_port, 
                           B(22) => q_6_1_22_port, B(21) => q_6_1_21_port, 
                           B(20) => q_6_1_20_port, B(19) => q_6_1_19_port, 
                           B(18) => q_6_1_18_port, B(17) => q_6_1_17_port, 
                           B(16) => q_6_1_16_port, B(15) => q_6_1_15_port, 
                           B(14) => q_6_1_14_port, B(13) => q_6_1_13_port, 
                           B(12) => q_6_1_12_port, B(11) => q_6_1_11_port, 
                           B(10) => q_6_1_10_port, B(9) => q_6_1_9_port, B(8) 
                           => q_6_1_8_port, B(7) => q_6_1_7_port, B(6) => 
                           q_6_1_6_port, B(5) => q_6_1_5_port, B(4) => 
                           q_6_1_4_port, B(3) => q_6_1_3_port, B(2) => B(3), 
                           B(1) => X_Logic0_port, B(0) => B(1), Cin => 
                           X_Logic0_port, S(63) => n_2062, S(62) => n_2063, 
                           S(61) => n_2064, S(60) => n_2065, S(59) => n_2066, 
                           S(58) => n_2067, S(57) => n_2068, S(56) => n_2069, 
                           S(55) => n_2070, S(54) => n_2071, S(53) => n_2072, 
                           S(52) => n_2073, S(51) => n_2074, S(50) => n_2075, 
                           S(49) => n_2076, S(48) => n_2077, S(47) => C(47), 
                           S(46) => C(46), S(45) => C(45), S(44) => C(44), 
                           S(43) => C(43), S(42) => C(42), S(41) => C(41), 
                           S(40) => C(40), S(39) => C(39), S(38) => C(38), 
                           S(37) => C(37), S(36) => C(36), S(35) => C(35), 
                           S(34) => C(34), S(33) => C(33), S(32) => C(32), 
                           S(31) => C(31), S(30) => C(30), S(29) => C(29), 
                           S(28) => C(28), S(27) => C(27), S(26) => C(26), 
                           S(25) => C(25), S(24) => C(24), S(23) => C(23), 
                           S(22) => C(22), S(21) => n_2078, S(20) => n_2079, 
                           S(19) => n_2080, S(18) => n_2081, S(17) => n_2082, 
                           S(16) => n_2083, S(15) => n_2084, S(14) => n_2085, 
                           S(13) => n_2086, S(12) => n_2087, S(11) => n_2088, 
                           S(10) => n_2089, S(9) => n_2090, S(8) => n_2091, 
                           S(7) => n_2092, S(6) => n_2093, S(5) => n_2094, S(4)
                           => n_2095, S(3) => n_2096, S(2) => n_2097, S(1) => 
                           n_2098, S(0) => n_2099, Cout => n_2100, clk => clk);
   U3 : BUF_X2 port map( A => A(23), Z => n381);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity UnpackFP_1 is

   port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector 
         (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, isNaN,
         isINF, isZ, isDN : out std_logic);

end UnpackFP_1;

architecture SYN_UnpackFP of UnpackFP_1 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N13, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13_port, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n_2101, 
      n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108 : std_logic;

begin
   SIG <= ( n_2101, n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, N13
      , FP(22), FP(21), FP(20), FP(19), FP(18), FP(17), FP(16), FP(15), FP(14),
      FP(13), FP(12), FP(11), FP(10), FP(9), FP(8), FP(7), FP(6), FP(5), FP(4),
      FP(3), FP(2), FP(1), FP(0) );
   EXP <= ( FP(30), FP(29), FP(28), FP(27), FP(26), FP(25), FP(24), FP(23) );
   SIGN <= FP(31);
   
   U2 : NAND4_X1 port map( A1 => n24, A2 => n23, A3 => n22, A4 => n21, ZN => 
                           n35);
   U3 : NOR2_X1 port map( A1 => FP(0), A2 => FP(1), ZN => n24);
   U4 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => n22);
   U5 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U6 : NOR2_X1 port map( A1 => FP(10), A2 => FP(9), ZN => n3);
   U7 : INV_X1 port map( A => FP(19), ZN => n17);
   U8 : INV_X1 port map( A => FP(20), ZN => n16);
   U9 : NOR2_X1 port map( A1 => FP(18), A2 => FP(17), ZN => n18);
   U10 : INV_X1 port map( A => FP(13), ZN => n12);
   U11 : INV_X1 port map( A => FP(14), ZN => n11);
   U12 : NOR2_X1 port map( A1 => FP(12), A2 => FP(11), ZN => n13_port);
   U13 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n23);
   U14 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n9);
   U15 : NAND4_X1 port map( A1 => n6, A2 => n5, A3 => n4, A4 => n3, ZN => n10);
   U16 : INV_X1 port map( A => FP(4), ZN => n7);
   U17 : NOR2_X1 port map( A1 => FP(3), A2 => FP(2), ZN => n8);
   U18 : NOR2_X1 port map( A1 => FP(5), A2 => FP(6), ZN => n6);
   U19 : OR2_X1 port map( A1 => FP(22), A2 => FP(21), ZN => n19);
   U20 : OR2_X1 port map( A1 => FP(16), A2 => FP(15), ZN => n14);
   U21 : INV_X1 port map( A => FP(8), ZN => n4);
   U22 : INV_X1 port map( A => FP(7), ZN => n5);
   U26 : NAND3_X1 port map( A1 => n13_port, A2 => n12, A3 => n11, ZN => n15);
   U27 : NAND3_X1 port map( A1 => n18, A2 => n17, A3 => n16, ZN => n20);
   U28 : INV_X1 port map( A => n35, ZN => n37);
   U30 : NOR2_X1 port map( A1 => N13, A2 => n35, ZN => isZ);
   U31 : INV_X1 port map( A => FP(28), ZN => n28);
   U32 : INV_X1 port map( A => FP(27), ZN => n27);
   U33 : INV_X1 port map( A => FP(30), ZN => n26);
   U34 : INV_X1 port map( A => FP(29), ZN => n25);
   U35 : NOR4_X1 port map( A1 => n28, A2 => n27, A3 => n26, A4 => n25, ZN => 
                           n34);
   U36 : INV_X1 port map( A => FP(24), ZN => n32);
   U37 : INV_X1 port map( A => FP(23), ZN => n31);
   U38 : INV_X1 port map( A => FP(26), ZN => n30);
   U39 : INV_X1 port map( A => FP(25), ZN => n29);
   U40 : NOR4_X1 port map( A1 => n32, A2 => n31, A3 => n30, A4 => n29, ZN => 
                           n33);
   U41 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => n36);
   U42 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => isINF);
   U43 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => isNaN);
   U23 : NAND2_X2 port map( A1 => n2, A2 => n1, ZN => N13);
   U24 : NOR2_X1 port map( A1 => FP(29), A2 => FP(30), ZN => n38);
   U25 : AND2_X1 port map( A1 => n39, A2 => n38, ZN => n2);
   U29 : NOR2_X1 port map( A1 => FP(27), A2 => FP(28), ZN => n39);
   U44 : NOR2_X1 port map( A1 => FP(25), A2 => FP(26), ZN => n40);
   U45 : AND2_X1 port map( A1 => n41, A2 => n40, ZN => n1);
   U46 : NOR2_X1 port map( A1 => FP(23), A2 => FP(24), ZN => n41);

end SYN_UnpackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity UnpackFP_0 is

   port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector 
         (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, isNaN,
         isINF, isZ, isDN : out std_logic);

end UnpackFP_0;

architecture SYN_UnpackFP of UnpackFP_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N13, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13_port, n14
      , n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, 
      n29, n30, n31, n32, n33, n34, n35, n36, n37, n_2110, n_2111, n_2112, 
      n_2113, n_2114, n_2115, n_2116, n_2117 : std_logic;

begin
   SIG <= ( n_2110, n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, N13
      , FP(22), FP(21), FP(20), FP(19), FP(18), FP(17), FP(16), FP(15), FP(14),
      FP(13), FP(12), FP(11), FP(10), FP(9), FP(8), FP(7), FP(6), FP(5), FP(4),
      FP(3), FP(2), FP(1), FP(0) );
   EXP <= ( FP(30), FP(29), FP(28), FP(27), FP(26), FP(25), FP(24), FP(23) );
   SIGN <= FP(31);
   
   U2 : NAND4_X1 port map( A1 => n24, A2 => n23, A3 => n22, A4 => n21, ZN => 
                           n35);
   U3 : NOR2_X1 port map( A1 => FP(0), A2 => FP(1), ZN => n24);
   U4 : NOR2_X1 port map( A1 => n15, A2 => n14, ZN => n22);
   U5 : NOR2_X1 port map( A1 => n20, A2 => n19, ZN => n21);
   U6 : NOR2_X1 port map( A1 => FP(10), A2 => FP(9), ZN => n3);
   U7 : INV_X1 port map( A => FP(19), ZN => n17);
   U8 : INV_X1 port map( A => FP(20), ZN => n16);
   U9 : NOR2_X1 port map( A1 => FP(18), A2 => FP(17), ZN => n18);
   U10 : INV_X1 port map( A => FP(13), ZN => n12);
   U11 : INV_X1 port map( A => FP(14), ZN => n11);
   U12 : NOR2_X1 port map( A1 => FP(12), A2 => FP(11), ZN => n13_port);
   U13 : NOR2_X1 port map( A1 => n10, A2 => n9, ZN => n23);
   U14 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => n9);
   U15 : NAND4_X1 port map( A1 => n6, A2 => n5, A3 => n4, A4 => n3, ZN => n10);
   U16 : INV_X1 port map( A => FP(4), ZN => n7);
   U17 : NOR2_X1 port map( A1 => FP(3), A2 => FP(2), ZN => n8);
   U18 : NOR2_X1 port map( A1 => FP(5), A2 => FP(6), ZN => n6);
   U19 : OR2_X1 port map( A1 => FP(22), A2 => FP(21), ZN => n19);
   U20 : OR2_X1 port map( A1 => FP(16), A2 => FP(15), ZN => n14);
   U21 : INV_X1 port map( A => FP(8), ZN => n4);
   U22 : INV_X1 port map( A => FP(7), ZN => n5);
   U23 : NOR4_X1 port map( A1 => FP(27), A2 => FP(28), A3 => FP(29), A4 => 
                           FP(30), ZN => n2);
   U26 : NAND3_X1 port map( A1 => n13_port, A2 => n12, A3 => n11, ZN => n15);
   U27 : NAND3_X1 port map( A1 => n18, A2 => n17, A3 => n16, ZN => n20);
   U28 : INV_X1 port map( A => n35, ZN => n37);
   U30 : NOR2_X1 port map( A1 => N13, A2 => n35, ZN => isZ);
   U31 : INV_X1 port map( A => FP(28), ZN => n28);
   U32 : INV_X1 port map( A => FP(27), ZN => n27);
   U33 : INV_X1 port map( A => FP(30), ZN => n26);
   U34 : INV_X1 port map( A => FP(29), ZN => n25);
   U35 : NOR4_X1 port map( A1 => n28, A2 => n27, A3 => n26, A4 => n25, ZN => 
                           n34);
   U36 : INV_X1 port map( A => FP(24), ZN => n32);
   U37 : INV_X1 port map( A => FP(23), ZN => n31);
   U38 : INV_X1 port map( A => FP(26), ZN => n30);
   U39 : INV_X1 port map( A => FP(25), ZN => n29);
   U40 : NOR4_X1 port map( A1 => n32, A2 => n31, A3 => n30, A4 => n29, ZN => 
                           n33);
   U41 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => n36);
   U42 : NOR2_X1 port map( A1 => n36, A2 => n35, ZN => isINF);
   U43 : NOR2_X1 port map( A1 => n37, A2 => n36, ZN => isNaN);
   U24 : NOR4_X1 port map( A1 => FP(23), A2 => FP(24), A3 => FP(25), A4 => 
                           FP(26), ZN => n1);
   U25 : NAND2_X1 port map( A1 => n2, A2 => n1, ZN => N13);

end SYN_UnpackFP;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage4 is

   port( EXP_neg : in std_logic;  EXP_out_round : in std_logic_vector (7 downto
         0);  EXP_pos, SIGN_out : in std_logic;  SIG_out_round : in 
         std_logic_vector (27 downto 0);  clk, isINF_tab, isNaN, isZ_tab : in 
         std_logic;  FP_Z : out std_logic_vector (31 downto 0));

end FPmul_stage4;

architecture SYN_struct of FPmul_stage4 is

   component PackFP
      port( SIGN : in std_logic;  EXP : in std_logic_vector (7 downto 0);  SIG 
            : in std_logic_vector (22 downto 0);  isNaN, isINF, isZ : in 
            std_logic;  FP : out std_logic_vector (31 downto 0);  clk : in 
            std_logic);
   end component;
   
   component FPnormalize_SIG_width28_1
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
            std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SIG_out_norm2_26_port, SIG_out_22_port, SIG_out_21_port, 
      SIG_out_20_port, SIG_out_19_port, SIG_out_18_port, SIG_out_17_port, 
      SIG_out_16_port, SIG_out_15_port, SIG_out_14_port, SIG_out_13_port, 
      SIG_out_12_port, SIG_out_11_port, SIG_out_10_port, SIG_out_9_port, 
      SIG_out_8_port, SIG_out_7_port, SIG_out_6_port, SIG_out_5_port, 
      SIG_out_4_port, SIG_out_3_port, SIG_out_2_port, SIG_out_1_port, 
      SIG_out_0_port, EXP_out_7_port, EXP_out_5_port, EXP_out_4_port, 
      EXP_out_3_port, EXP_out_2_port, EXP_out_1_port, EXP_out_0_port, isINF, n1
      , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n24,
      n25, n26, n32, n33, n47, n49, n116, n117, n118, n122, n123, n124, n125, 
      n144, n145, n146, n147, n148, n149, n150, n151, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, 
      n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, 
      n_2138, n_2139, n_2140, n_2141, n_2142, n_2143 : std_logic;

begin
   
   U6 : INV_X1 port map( A => EXP_out_0_port, ZN => n24);
   U7 : INV_X1 port map( A => EXP_out_2_port, ZN => n25);
   U9 : INV_X1 port map( A => isINF_tab, ZN => n49);
   U10 : INV_X1 port map( A => EXP_pos, ZN => n47);
   U11 : NOR2_X1 port map( A1 => n25, A2 => n24, ZN => n26);
   U12 : INV_X1 port map( A => SIG_out_5_port, ZN => n4);
   U13 : INV_X1 port map( A => SIG_out_4_port, ZN => n3);
   U14 : INV_X1 port map( A => SIG_out_3_port, ZN => n2);
   U15 : NOR3_X1 port map( A1 => n159, A2 => n160, A3 => n161, ZN => n1);
   U17 : INV_X1 port map( A => SIG_out_11_port, ZN => n8);
   U18 : INV_X1 port map( A => SIG_out_10_port, ZN => n7);
   U19 : INV_X1 port map( A => SIG_out_9_port, ZN => n6);
   U22 : INV_X1 port map( A => SIG_out_17_port, ZN => n12);
   U23 : INV_X1 port map( A => SIG_out_16_port, ZN => n11);
   U24 : INV_X1 port map( A => SIG_out_15_port, ZN => n10);
   U25 : NOR3_X1 port map( A1 => SIG_out_14_port, A2 => SIG_out_13_port, A3 => 
                           SIG_out_12_port, ZN => n9);
   U27 : INV_X1 port map( A => SIG_out_20_port, ZN => n16);
   U28 : INV_X1 port map( A => SIG_out_19_port, ZN => n15);
   U29 : INV_X1 port map( A => SIG_out_18_port, ZN => n14);
   U30 : NOR3_X1 port map( A1 => SIG_out_21_port, A2 => SIG_out_22_port, A3 => 
                           SIG_out_norm2_26_port, ZN => n13);
   n116 <= '0';
   n117 <= '0';
   n118 <= '0';
   U31 : AND4_X1 port map( A1 => n4, A2 => n3, A3 => n2, A4 => n1, ZN => n122);
   U32 : AND4_X1 port map( A1 => n5, A2 => n7, A3 => n6, A4 => n8, ZN => n123);
   U37 : AND4_X1 port map( A1 => n9, A2 => n11, A3 => n10, A4 => n12, ZN => 
                           n124);
   U38 : AND4_X1 port map( A1 => n13, A2 => n15, A3 => n14, A4 => n16, ZN => 
                           n125);
   MY_CLK_r_REG206_S4 : DFF_X1 port map( D => SIG_out_2_port, CK => clk, Q => 
                           n161, QN => n_2122);
   MY_CLK_r_REG207_S4 : DFF_X1 port map( D => SIG_out_1_port, CK => clk, Q => 
                           n160, QN => n_2123);
   MY_CLK_r_REG208_S4 : DFF_X1 port map( D => SIG_out_0_port, CK => clk, Q => 
                           n159, QN => n_2124);
   MY_CLK_r_REG196_S1 : DFF_X1 port map( D => n49, CK => clk, Q => n158, QN => 
                           n_2125);
   MY_CLK_r_REG197_S2 : DFF_X1 port map( D => n158, CK => clk, Q => n157, QN =>
                           n_2126);
   MY_CLK_r_REG198_S3 : DFF_X1 port map( D => n157, CK => clk, Q => n156, QN =>
                           n_2127);
   MY_CLK_r_REG199_S4 : DFF_X1 port map( D => n156, CK => clk, Q => n155, QN =>
                           n_2128);
   MY_CLK_r_REG383_S2 : DFF_X1 port map( D => n47, CK => clk, Q => n154, QN => 
                           n_2129);
   MY_CLK_r_REG384_S3 : DFF_X1 port map( D => n154, CK => clk, Q => n153, QN =>
                           n_2130);
   MY_CLK_r_REG385_S4 : DFF_X1 port map( D => n153, CK => clk, Q => n_2131, QN 
                           => n181);
   MY_CLK_r_REG379_S1 : DFF_X1 port map( D => EXP_neg, CK => clk, Q => n151, QN
                           => n_2132);
   MY_CLK_r_REG380_S2 : DFF_X1 port map( D => n151, CK => clk, Q => n150, QN =>
                           n_2133);
   MY_CLK_r_REG381_S3 : DFF_X1 port map( D => n150, CK => clk, Q => n149, QN =>
                           n_2134);
   MY_CLK_r_REG382_S4 : DFF_X1 port map( D => n149, CK => clk, Q => n148, QN =>
                           n_2135);
   MY_CLK_r_REG192_S1 : DFF_X1 port map( D => isZ_tab, CK => clk, Q => n147, QN
                           => n_2136);
   MY_CLK_r_REG193_S2 : DFF_X1 port map( D => n147, CK => clk, Q => n146, QN =>
                           n_2137);
   MY_CLK_r_REG194_S3 : DFF_X1 port map( D => n146, CK => clk, Q => n145, QN =>
                           n_2138);
   MY_CLK_r_REG195_S4 : DFF_X1 port map( D => n145, CK => clk, Q => n144, QN =>
                           n_2139);
   U3 : AND2_X1 port map( A1 => n180, A2 => EXP_out_5_port, ZN => n186);
   U4 : AND2_X1 port map( A1 => EXP_out_3_port, A2 => EXP_out_4_port, ZN => 
                           n185);
   U5 : AOI21_X1 port map( B1 => n32, B2 => n155, A => n33, ZN => isINF);
   U8 : NAND2_X1 port map( A1 => n187, A2 => n188, ZN => n33);
   U20 : NAND2_X1 port map( A1 => n183, A2 => n182, ZN => n32);
   U21 : OR2_X1 port map( A1 => EXP_out_7_port, A2 => n181, ZN => n182);
   U26 : NAND2_X1 port map( A1 => n184, A2 => EXP_out_7_port, ZN => n183);
   U33 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => EXP_out_1_port, A4 =>
                           n26, ZN => n184);
   U34 : NAND4_X1 port map( A1 => n124, A2 => n123, A3 => n125, A4 => n122, ZN 
                           => n188);
   U35 : AOI21_X1 port map( B1 => EXP_out_7_port, B2 => n148, A => n144, ZN => 
                           n187);
   U36 : NOR3_X1 port map( A1 => SIG_out_8_port, A2 => SIG_out_6_port, A3 => 
                           SIG_out_7_port, ZN => n5);
   I1 : FPnormalize_SIG_width28_1 port map( SIG_in(27) => SIG_out_round(27), 
                           SIG_in(26) => SIG_out_round(26), SIG_in(25) => 
                           SIG_out_round(25), SIG_in(24) => SIG_out_round(24), 
                           SIG_in(23) => SIG_out_round(23), SIG_in(22) => 
                           SIG_out_round(22), SIG_in(21) => SIG_out_round(21), 
                           SIG_in(20) => SIG_out_round(20), SIG_in(19) => 
                           SIG_out_round(19), SIG_in(18) => SIG_out_round(18), 
                           SIG_in(17) => SIG_out_round(17), SIG_in(16) => 
                           SIG_out_round(16), SIG_in(15) => SIG_out_round(15), 
                           SIG_in(14) => SIG_out_round(14), SIG_in(13) => 
                           SIG_out_round(13), SIG_in(12) => SIG_out_round(12), 
                           SIG_in(11) => SIG_out_round(11), SIG_in(10) => 
                           SIG_out_round(10), SIG_in(9) => SIG_out_round(9), 
                           SIG_in(8) => SIG_out_round(8), SIG_in(7) => 
                           SIG_out_round(7), SIG_in(6) => SIG_out_round(6), 
                           SIG_in(5) => SIG_out_round(5), SIG_in(4) => 
                           SIG_out_round(4), SIG_in(3) => SIG_out_round(3), 
                           SIG_in(2) => n116, SIG_in(1) => n117, SIG_in(0) => 
                           n118, EXP_in(7) => EXP_out_round(7), EXP_in(6) => 
                           EXP_out_round(6), EXP_in(5) => EXP_out_round(5), 
                           EXP_in(4) => EXP_out_round(4), EXP_in(3) => 
                           EXP_out_round(3), EXP_in(2) => EXP_out_round(2), 
                           EXP_in(1) => EXP_out_round(1), EXP_in(0) => 
                           EXP_out_round(0), SIG_out(27) => n_2140, SIG_out(26)
                           => SIG_out_norm2_26_port, SIG_out(25) => 
                           SIG_out_22_port, SIG_out(24) => SIG_out_21_port, 
                           SIG_out(23) => SIG_out_20_port, SIG_out(22) => 
                           SIG_out_19_port, SIG_out(21) => SIG_out_18_port, 
                           SIG_out(20) => SIG_out_17_port, SIG_out(19) => 
                           SIG_out_16_port, SIG_out(18) => SIG_out_15_port, 
                           SIG_out(17) => SIG_out_14_port, SIG_out(16) => 
                           SIG_out_13_port, SIG_out(15) => SIG_out_12_port, 
                           SIG_out(14) => SIG_out_11_port, SIG_out(13) => 
                           SIG_out_10_port, SIG_out(12) => SIG_out_9_port, 
                           SIG_out(11) => SIG_out_8_port, SIG_out(10) => 
                           SIG_out_7_port, SIG_out(9) => SIG_out_6_port, 
                           SIG_out(8) => SIG_out_5_port, SIG_out(7) => 
                           SIG_out_4_port, SIG_out(6) => SIG_out_3_port, 
                           SIG_out(5) => SIG_out_2_port, SIG_out(4) => 
                           SIG_out_1_port, SIG_out(3) => SIG_out_0_port, 
                           SIG_out(2) => n_2141, SIG_out(1) => n_2142, 
                           SIG_out(0) => n_2143, EXP_out(7) => EXP_out_7_port, 
                           EXP_out(6) => n180, EXP_out(5) => EXP_out_5_port, 
                           EXP_out(4) => EXP_out_4_port, EXP_out(3) => 
                           EXP_out_3_port, EXP_out(2) => EXP_out_2_port, 
                           EXP_out(1) => EXP_out_1_port, EXP_out(0) => 
                           EXP_out_0_port, clk => clk);
   I3 : PackFP port map( SIGN => SIGN_out, EXP(7) => EXP_out_7_port, EXP(6) => 
                           n180, EXP(5) => EXP_out_5_port, EXP(4) => 
                           EXP_out_4_port, EXP(3) => EXP_out_3_port, EXP(2) => 
                           EXP_out_2_port, EXP(1) => EXP_out_1_port, EXP(0) => 
                           EXP_out_0_port, SIG(22) => SIG_out_22_port, SIG(21) 
                           => SIG_out_21_port, SIG(20) => SIG_out_20_port, 
                           SIG(19) => SIG_out_19_port, SIG(18) => 
                           SIG_out_18_port, SIG(17) => SIG_out_17_port, SIG(16)
                           => SIG_out_16_port, SIG(15) => SIG_out_15_port, 
                           SIG(14) => SIG_out_14_port, SIG(13) => 
                           SIG_out_13_port, SIG(12) => SIG_out_12_port, SIG(11)
                           => SIG_out_11_port, SIG(10) => SIG_out_10_port, 
                           SIG(9) => SIG_out_9_port, SIG(8) => SIG_out_8_port, 
                           SIG(7) => SIG_out_7_port, SIG(6) => SIG_out_6_port, 
                           SIG(5) => SIG_out_5_port, SIG(4) => SIG_out_4_port, 
                           SIG(3) => SIG_out_3_port, SIG(2) => n161, SIG(1) => 
                           n160, SIG(0) => n159, isNaN => isNaN, isINF => isINF
                           , isZ => n33, FP(31) => FP_Z(31), FP(30) => FP_Z(30)
                           , FP(29) => FP_Z(29), FP(28) => FP_Z(28), FP(27) => 
                           FP_Z(27), FP(26) => FP_Z(26), FP(25) => FP_Z(25), 
                           FP(24) => FP_Z(24), FP(23) => FP_Z(23), FP(22) => 
                           FP_Z(22), FP(21) => FP_Z(21), FP(20) => FP_Z(20), 
                           FP(19) => FP_Z(19), FP(18) => FP_Z(18), FP(17) => 
                           FP_Z(17), FP(16) => FP_Z(16), FP(15) => FP_Z(15), 
                           FP(14) => FP_Z(14), FP(13) => FP_Z(13), FP(12) => 
                           FP_Z(12), FP(11) => FP_Z(11), FP(10) => FP_Z(10), 
                           FP(9) => FP_Z(9), FP(8) => FP_Z(8), FP(7) => FP_Z(7)
                           , FP(6) => FP_Z(6), FP(5) => FP_Z(5), FP(4) => 
                           FP_Z(4), FP(3) => FP_Z(3), FP(2) => FP_Z(2), FP(1) 
                           => FP_Z(1), FP(0) => FP_Z(0), clk => clk);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage3 is

   port( EXP_in : in std_logic_vector (7 downto 0);  EXP_neg_stage2, 
         EXP_pos_stage2, SIGN_out_stage2 : in std_logic;  SIG_in : in 
         std_logic_vector (27 downto 0);  clk, isINF_stage2, isNaN_stage2, 
         isZ_tab_stage2 : in std_logic;  EXP_neg : out std_logic;  
         EXP_out_round : out std_logic_vector (7 downto 0);  EXP_pos, SIGN_out 
         : out std_logic;  SIG_out_round : out std_logic_vector (27 downto 0); 
         isINF_tab, isNaN, isZ_tab : out std_logic);

end FPmul_stage3;

architecture SYN_struct of FPmul_stage3 is

   component FPround_SIG_width28
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0));
   end component;
   
   component FPnormalize_SIG_width28_0
      port( SIG_in : in std_logic_vector (27 downto 0);  EXP_in : in 
            std_logic_vector (7 downto 0);  SIG_out : out std_logic_vector (27 
            downto 0);  EXP_out : out std_logic_vector (7 downto 0);  clk : in 
            std_logic);
   end component;
   
   signal SIG_out_norm_27_port, SIG_out_norm_26_port, SIG_out_norm_25_port, 
      SIG_out_norm_24_port, SIG_out_norm_23_port, SIG_out_norm_22_port, 
      SIG_out_norm_21_port, SIG_out_norm_20_port, SIG_out_norm_19_port, 
      SIG_out_norm_18_port, SIG_out_norm_17_port, SIG_out_norm_16_port, 
      SIG_out_norm_14_port, SIG_out_norm_13_port, SIG_out_norm_10_port, 
      SIG_out_norm_9_port, SIG_out_norm_8_port, SIG_out_norm_7_port, 
      SIG_out_norm_6_port, SIG_out_norm_5_port, SIG_out_norm_4_port, 
      SIG_out_norm_3_port, SIG_out_norm_2_port, EXP_out_norm_7_port, 
      EXP_out_norm_6_port, EXP_out_norm_5_port, EXP_out_norm_4_port, 
      EXP_out_norm_3_port, EXP_out_norm_2_port, EXP_out_norm_1_port, 
      EXP_out_norm_0_port, n79, n80, n81, n82, n83, n84, n85, n_2149, n_2150, 
      n_2151, n_2152, n_2153, n_2154 : std_logic;

begin
   EXP_neg <= EXP_neg_stage2;
   EXP_pos <= EXP_pos_stage2;
   SIGN_out <= SIGN_out_stage2;
   isINF_tab <= isINF_stage2;
   isNaN <= isNaN_stage2;
   isZ_tab <= isZ_tab_stage2;
   
   SIG_out_norm_27_port <= '0';
   n79 <= '0';
   n80 <= '0';
   n81 <= '0';
   n82 <= '0';
   I9 : FPnormalize_SIG_width28_0 port map( SIG_in(27) => SIG_in(27), 
                           SIG_in(26) => SIG_in(26), SIG_in(25) => SIG_in(25), 
                           SIG_in(24) => SIG_in(24), SIG_in(23) => SIG_in(23), 
                           SIG_in(22) => SIG_in(22), SIG_in(21) => SIG_in(21), 
                           SIG_in(20) => SIG_in(20), SIG_in(19) => SIG_in(19), 
                           SIG_in(18) => SIG_in(18), SIG_in(17) => SIG_in(17), 
                           SIG_in(16) => SIG_in(16), SIG_in(15) => SIG_in(15), 
                           SIG_in(14) => SIG_in(14), SIG_in(13) => SIG_in(13), 
                           SIG_in(12) => SIG_in(12), SIG_in(11) => SIG_in(11), 
                           SIG_in(10) => SIG_in(10), SIG_in(9) => SIG_in(9), 
                           SIG_in(8) => SIG_in(8), SIG_in(7) => SIG_in(7), 
                           SIG_in(6) => SIG_in(6), SIG_in(5) => SIG_in(5), 
                           SIG_in(4) => SIG_in(4), SIG_in(3) => SIG_in(3), 
                           SIG_in(2) => SIG_in(2), SIG_in(1) => n79, SIG_in(0) 
                           => n80, EXP_in(7) => EXP_in(7), EXP_in(6) => 
                           EXP_in(6), EXP_in(5) => EXP_in(5), EXP_in(4) => 
                           EXP_in(4), EXP_in(3) => EXP_in(3), EXP_in(2) => 
                           EXP_in(2), EXP_in(1) => EXP_in(1), EXP_in(0) => 
                           EXP_in(0), SIG_out(27) => n_2149, SIG_out(26) => 
                           SIG_out_norm_26_port, SIG_out(25) => 
                           SIG_out_norm_25_port, SIG_out(24) => 
                           SIG_out_norm_24_port, SIG_out(23) => 
                           SIG_out_norm_23_port, SIG_out(22) => 
                           SIG_out_norm_22_port, SIG_out(21) => 
                           SIG_out_norm_21_port, SIG_out(20) => 
                           SIG_out_norm_20_port, SIG_out(19) => 
                           SIG_out_norm_19_port, SIG_out(18) => 
                           SIG_out_norm_18_port, SIG_out(17) => 
                           SIG_out_norm_17_port, SIG_out(16) => 
                           SIG_out_norm_16_port, SIG_out(15) => n83, 
                           SIG_out(14) => SIG_out_norm_14_port, SIG_out(13) => 
                           SIG_out_norm_13_port, SIG_out(12) => n85, 
                           SIG_out(11) => n84, SIG_out(10) => 
                           SIG_out_norm_10_port, SIG_out(9) => 
                           SIG_out_norm_9_port, SIG_out(8) => 
                           SIG_out_norm_8_port, SIG_out(7) => 
                           SIG_out_norm_7_port, SIG_out(6) => 
                           SIG_out_norm_6_port, SIG_out(5) => 
                           SIG_out_norm_5_port, SIG_out(4) => 
                           SIG_out_norm_4_port, SIG_out(3) => 
                           SIG_out_norm_3_port, SIG_out(2) => 
                           SIG_out_norm_2_port, SIG_out(1) => n_2150, 
                           SIG_out(0) => n_2151, EXP_out(7) => 
                           EXP_out_norm_7_port, EXP_out(6) => 
                           EXP_out_norm_6_port, EXP_out(5) => 
                           EXP_out_norm_5_port, EXP_out(4) => 
                           EXP_out_norm_4_port, EXP_out(3) => 
                           EXP_out_norm_3_port, EXP_out(2) => 
                           EXP_out_norm_2_port, EXP_out(1) => 
                           EXP_out_norm_1_port, EXP_out(0) => 
                           EXP_out_norm_0_port, clk => clk);
   I11 : FPround_SIG_width28 port map( SIG_in(27) => SIG_out_norm_27_port, 
                           SIG_in(26) => SIG_out_norm_26_port, SIG_in(25) => 
                           SIG_out_norm_25_port, SIG_in(24) => 
                           SIG_out_norm_24_port, SIG_in(23) => 
                           SIG_out_norm_23_port, SIG_in(22) => 
                           SIG_out_norm_22_port, SIG_in(21) => 
                           SIG_out_norm_21_port, SIG_in(20) => 
                           SIG_out_norm_20_port, SIG_in(19) => 
                           SIG_out_norm_19_port, SIG_in(18) => 
                           SIG_out_norm_18_port, SIG_in(17) => 
                           SIG_out_norm_17_port, SIG_in(16) => 
                           SIG_out_norm_16_port, SIG_in(15) => n83, SIG_in(14) 
                           => SIG_out_norm_14_port, SIG_in(13) => 
                           SIG_out_norm_13_port, SIG_in(12) => n85, SIG_in(11) 
                           => n84, SIG_in(10) => SIG_out_norm_10_port, 
                           SIG_in(9) => SIG_out_norm_9_port, SIG_in(8) => 
                           SIG_out_norm_8_port, SIG_in(7) => 
                           SIG_out_norm_7_port, SIG_in(6) => 
                           SIG_out_norm_6_port, SIG_in(5) => 
                           SIG_out_norm_5_port, SIG_in(4) => 
                           SIG_out_norm_4_port, SIG_in(3) => 
                           SIG_out_norm_3_port, SIG_in(2) => 
                           SIG_out_norm_2_port, SIG_in(1) => n81, SIG_in(0) => 
                           n82, EXP_in(7) => EXP_out_norm_7_port, EXP_in(6) => 
                           EXP_out_norm_6_port, EXP_in(5) => 
                           EXP_out_norm_5_port, EXP_in(4) => 
                           EXP_out_norm_4_port, EXP_in(3) => 
                           EXP_out_norm_3_port, EXP_in(2) => 
                           EXP_out_norm_2_port, EXP_in(1) => 
                           EXP_out_norm_1_port, EXP_in(0) => 
                           EXP_out_norm_0_port, SIG_out(27) => 
                           SIG_out_round(27), SIG_out(26) => SIG_out_round(26),
                           SIG_out(25) => SIG_out_round(25), SIG_out(24) => 
                           SIG_out_round(24), SIG_out(23) => SIG_out_round(23),
                           SIG_out(22) => SIG_out_round(22), SIG_out(21) => 
                           SIG_out_round(21), SIG_out(20) => SIG_out_round(20),
                           SIG_out(19) => SIG_out_round(19), SIG_out(18) => 
                           SIG_out_round(18), SIG_out(17) => SIG_out_round(17),
                           SIG_out(16) => SIG_out_round(16), SIG_out(15) => 
                           SIG_out_round(15), SIG_out(14) => SIG_out_round(14),
                           SIG_out(13) => SIG_out_round(13), SIG_out(12) => 
                           SIG_out_round(12), SIG_out(11) => SIG_out_round(11),
                           SIG_out(10) => SIG_out_round(10), SIG_out(9) => 
                           SIG_out_round(9), SIG_out(8) => SIG_out_round(8), 
                           SIG_out(7) => SIG_out_round(7), SIG_out(6) => 
                           SIG_out_round(6), SIG_out(5) => SIG_out_round(5), 
                           SIG_out(4) => SIG_out_round(4), SIG_out(3) => 
                           SIG_out_round(3), SIG_out(2) => n_2152, SIG_out(1) 
                           => n_2153, SIG_out(0) => n_2154, EXP_out(7) => 
                           EXP_out_round(7), EXP_out(6) => EXP_out_round(6), 
                           EXP_out(5) => EXP_out_round(5), EXP_out(4) => 
                           EXP_out_round(4), EXP_out(3) => EXP_out_round(3), 
                           EXP_out(2) => EXP_out_round(2), EXP_out(1) => 
                           EXP_out_round(1), EXP_out(0) => EXP_out_round(0));

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage2 is

   port( A_EXP : in std_logic_vector (7 downto 0);  A_SIG : in std_logic_vector
         (31 downto 0);  B_EXP : in std_logic_vector (7 downto 0);  B_SIG : in 
         std_logic_vector (31 downto 0);  SIGN_out_stage1, clk, isINF_stage1, 
         isNaN_stage1, isZ_tab_stage1 : in std_logic;  EXP_in : out 
         std_logic_vector (7 downto 0);  EXP_neg_stage2, EXP_pos_stage2, 
         SIGN_out_stage2 : out std_logic;  SIG_in : out std_logic_vector (27 
         downto 0);  isINF_stage2, isNaN_stage2, isZ_tab_stage2 : out std_logic
         );

end FPmul_stage2;

architecture SYN_struct of FPmul_stage2 is

   component MBE
      port( A, B : in std_logic_vector (31 downto 0);  C : out std_logic_vector
            (63 downto 0);  clk : in std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
      n105, n106, n107, mw_I4sum_7_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, 
      n10, n110, n111, add_1_root_add_131_2_n6, add_1_root_add_131_2_n5, 
      add_1_root_add_131_2_n4, add_1_root_add_131_2_carry_1_port, 
      add_1_root_add_131_2_carry_2_port, add_1_root_add_131_2_carry_3_port, 
      add_1_root_add_131_2_carry_4_port, add_1_root_add_131_2_carry_5_port, 
      add_1_root_add_131_2_carry_6_port, add_1_root_add_131_2_carry_7_port, 
      n_2173, n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, 
      n_2182, n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, 
      n_2191, n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, 
      n_2200, n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, 
      n_2209, n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216 : 
      std_logic;

begin
   SIGN_out_stage2 <= SIGN_out_stage1;
   isINF_stage2 <= isINF_stage1;
   isNaN_stage2 <= isNaN_stage1;
   isZ_tab_stage2 <= isZ_tab_stage1;
   
   U3 : AND2_X1 port map( A1 => n111, A2 => n110, ZN => EXP_pos_stage2);
   U4 : NAND4_X1 port map( A1 => B_EXP(5), A2 => B_EXP(6), A3 => B_EXP(3), A4 
                           => B_EXP(4), ZN => n4);
   U5 : INV_X1 port map( A => B_EXP(0), ZN => n3);
   U6 : INV_X1 port map( A => B_EXP(2), ZN => n2);
   U7 : INV_X1 port map( A => B_EXP(1), ZN => n1);
   U8 : NOR4_X1 port map( A1 => n4, A2 => n3, A3 => n2, A4 => n1, ZN => n10);
   U9 : NAND4_X1 port map( A1 => A_EXP(5), A2 => A_EXP(6), A3 => A_EXP(3), A4 
                           => A_EXP(4), ZN => n8);
   U10 : INV_X1 port map( A => A_EXP(0), ZN => n7);
   U11 : INV_X1 port map( A => A_EXP(2), ZN => n6);
   U12 : INV_X1 port map( A => A_EXP(1), ZN => n5);
   U13 : NOR4_X1 port map( A1 => n8, A2 => n7, A3 => n6, A4 => n5, ZN => n9);
   U14 : NOR4_X1 port map( A1 => B_EXP(7), A2 => A_EXP(7), A3 => n10, A4 => n9,
                           ZN => EXP_neg_stage2);
   U15 : INV_X1 port map( A => mw_I4sum_7_port, ZN => EXP_in(7));
   n107 <= '0';
   n106 <= '0';
   n105 <= '0';
   n104 <= '0';
   n103 <= '0';
   n102 <= '0';
   n101 <= '0';
   n100 <= '0';
   n99 <= '0';
   n98 <= '0';
   n97 <= '0';
   n96 <= '0';
   n95 <= '0';
   n94 <= '0';
   n93 <= '0';
   n92 <= '0';
   MY_CLK_r_REG378_S1 : DFF_X1 port map( D => A_EXP(7), CK => clk, Q => n111, 
                           QN => n_2173);
   MY_CLK_r_REG639_S1 : DFF_X1 port map( D => B_EXP(7), CK => clk, Q => n110, 
                           QN => n_2174);
   add_1_root_add_131_2_MY_CLK_r_REG391_S1 : DFF_X1 port map( D => 
                           add_1_root_add_131_2_carry_6_port, CK => clk, Q => 
                           add_1_root_add_131_2_n4, QN => n_2175);
   add_1_root_add_131_2_MY_CLK_r_REG640_S1 : DFF_X1 port map( D => B_EXP(6), CK
                           => clk, Q => add_1_root_add_131_2_n5, QN => n_2176);
   add_1_root_add_131_2_MY_CLK_r_REG388_S1 : DFF_X1 port map( D => A_EXP(6), CK
                           => clk, Q => add_1_root_add_131_2_n6, QN => n_2177);
   add_1_root_add_131_2_U2 : XNOR2_X1 port map( A => B_EXP(0), B => A_EXP(0), 
                           ZN => EXP_in(0));
   add_1_root_add_131_2_U1 : OR2_X1 port map( A1 => B_EXP(0), A2 => A_EXP(0), 
                           ZN => add_1_root_add_131_2_carry_1_port);
   add_1_root_add_131_2_U1_1 : FA_X1 port map( A => A_EXP(1), B => B_EXP(1), CI
                           => add_1_root_add_131_2_carry_1_port, CO => 
                           add_1_root_add_131_2_carry_2_port, S => EXP_in(1));
   add_1_root_add_131_2_U1_2 : FA_X1 port map( A => A_EXP(2), B => B_EXP(2), CI
                           => add_1_root_add_131_2_carry_2_port, CO => 
                           add_1_root_add_131_2_carry_3_port, S => EXP_in(2));
   add_1_root_add_131_2_U1_3 : FA_X1 port map( A => A_EXP(3), B => B_EXP(3), CI
                           => add_1_root_add_131_2_carry_3_port, CO => 
                           add_1_root_add_131_2_carry_4_port, S => EXP_in(3));
   add_1_root_add_131_2_U1_4 : FA_X1 port map( A => A_EXP(4), B => B_EXP(4), CI
                           => add_1_root_add_131_2_carry_4_port, CO => 
                           add_1_root_add_131_2_carry_5_port, S => EXP_in(4));
   add_1_root_add_131_2_U1_5 : FA_X1 port map( A => A_EXP(5), B => B_EXP(5), CI
                           => add_1_root_add_131_2_carry_5_port, CO => 
                           add_1_root_add_131_2_carry_6_port, S => EXP_in(5));
   add_1_root_add_131_2_U1_6 : FA_X1 port map( A => add_1_root_add_131_2_n6, B 
                           => add_1_root_add_131_2_n5, CI => 
                           add_1_root_add_131_2_n4, CO => 
                           add_1_root_add_131_2_carry_7_port, S => EXP_in(6));
   add_1_root_add_131_2_U1_7 : FA_X1 port map( A => n111, B => n110, CI => 
                           add_1_root_add_131_2_carry_7_port, CO => n_2178, S 
                           => mw_I4sum_7_port);
   MBE_SIG : MBE port map( A(31) => n92, A(30) => n93, A(29) => n94, A(28) => 
                           n95, A(27) => n96, A(26) => n97, A(25) => n98, A(24)
                           => n99, A(23) => A_SIG(23), A(22) => A_SIG(22), 
                           A(21) => A_SIG(21), A(20) => A_SIG(20), A(19) => 
                           A_SIG(19), A(18) => A_SIG(18), A(17) => A_SIG(17), 
                           A(16) => A_SIG(16), A(15) => A_SIG(15), A(14) => 
                           A_SIG(14), A(13) => A_SIG(13), A(12) => A_SIG(12), 
                           A(11) => A_SIG(11), A(10) => A_SIG(10), A(9) => 
                           A_SIG(9), A(8) => A_SIG(8), A(7) => A_SIG(7), A(6) 
                           => A_SIG(6), A(5) => A_SIG(5), A(4) => A_SIG(4), 
                           A(3) => A_SIG(3), A(2) => A_SIG(2), A(1) => A_SIG(1)
                           , A(0) => A_SIG(0), B(31) => n100, B(30) => n101, 
                           B(29) => n102, B(28) => n103, B(27) => n104, B(26) 
                           => n105, B(25) => n106, B(24) => n107, B(23) => 
                           B_SIG(23), B(22) => B_SIG(22), B(21) => B_SIG(21), 
                           B(20) => B_SIG(20), B(19) => B_SIG(19), B(18) => 
                           B_SIG(18), B(17) => B_SIG(17), B(16) => B_SIG(16), 
                           B(15) => B_SIG(15), B(14) => B_SIG(14), B(13) => 
                           B_SIG(13), B(12) => B_SIG(12), B(11) => B_SIG(11), 
                           B(10) => B_SIG(10), B(9) => B_SIG(9), B(8) => 
                           B_SIG(8), B(7) => B_SIG(7), B(6) => B_SIG(6), B(5) 
                           => B_SIG(5), B(4) => B_SIG(4), B(3) => B_SIG(3), 
                           B(2) => B_SIG(2), B(1) => B_SIG(1), B(0) => B_SIG(0)
                           , C(63) => n_2179, C(62) => n_2180, C(61) => n_2181,
                           C(60) => n_2182, C(59) => n_2183, C(58) => n_2184, 
                           C(57) => n_2185, C(56) => n_2186, C(55) => n_2187, 
                           C(54) => n_2188, C(53) => n_2189, C(52) => n_2190, 
                           C(51) => n_2191, C(50) => n_2192, C(49) => n_2193, 
                           C(48) => n_2194, C(47) => SIG_in(27), C(46) => 
                           SIG_in(26), C(45) => SIG_in(25), C(44) => SIG_in(24)
                           , C(43) => SIG_in(23), C(42) => SIG_in(22), C(41) =>
                           SIG_in(21), C(40) => SIG_in(20), C(39) => SIG_in(19)
                           , C(38) => SIG_in(18), C(37) => SIG_in(17), C(36) =>
                           SIG_in(16), C(35) => SIG_in(15), C(34) => SIG_in(14)
                           , C(33) => SIG_in(13), C(32) => SIG_in(12), C(31) =>
                           SIG_in(11), C(30) => SIG_in(10), C(29) => SIG_in(9),
                           C(28) => SIG_in(8), C(27) => SIG_in(7), C(26) => 
                           SIG_in(6), C(25) => SIG_in(5), C(24) => SIG_in(4), 
                           C(23) => SIG_in(3), C(22) => SIG_in(2), C(21) => 
                           n_2195, C(20) => n_2196, C(19) => n_2197, C(18) => 
                           n_2198, C(17) => n_2199, C(16) => n_2200, C(15) => 
                           n_2201, C(14) => n_2202, C(13) => n_2203, C(12) => 
                           n_2204, C(11) => n_2205, C(10) => n_2206, C(9) => 
                           n_2207, C(8) => n_2208, C(7) => n_2209, C(6) => 
                           n_2210, C(5) => n_2211, C(4) => n_2212, C(3) => 
                           n_2213, C(2) => n_2214, C(1) => n_2215, C(0) => 
                           n_2216, clk => clk);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul_stage1 is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         A_EXP : out std_logic_vector (7 downto 0);  A_SIG : out 
         std_logic_vector (31 downto 0);  B_EXP : out std_logic_vector (7 
         downto 0);  B_SIG : out std_logic_vector (31 downto 0);  
         SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : out 
         std_logic);

end FPmul_stage1;

architecture SYN_struct of FPmul_stage1 is

   component UnpackFP_1
      port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector
            (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, 
            isNaN, isINF, isZ, isDN : out std_logic);
   end component;
   
   component UnpackFP_0
      port( FP : in std_logic_vector (31 downto 0);  SIG : out std_logic_vector
            (31 downto 0);  EXP : out std_logic_vector (7 downto 0);  SIGN, 
            isNaN, isINF, isZ, isDN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal A_isINF, A_isNaN, A_isZ, B_isINF, B_isNaN, B_isZ, A_SIGN, B_SIGN, n18
      , n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n_2233, n_2234, 
      n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, 
      n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250 : std_logic;

begin
   
   U25 : INV_X1 port map( A => B_isZ, ZN => n20);
   U26 : INV_X1 port map( A => A_isZ, ZN => n22);
   U27 : OR2_X1 port map( A1 => B_isNaN, A2 => A_isNaN, ZN => n21);
   U28 : INV_X1 port map( A => n21, ZN => n18);
   U29 : INV_X1 port map( A => A_isINF, ZN => n25);
   U30 : NAND2_X1 port map( A1 => n18, A2 => n25, ZN => n19);
   U31 : AOI211_X1 port map( C1 => n20, C2 => n22, A => n19, B => B_isINF, ZN 
                           => isZ_tab_stage1);
   U32 : NAND2_X1 port map( A1 => B_isZ, A2 => A_isINF, ZN => n26);
   U33 : NAND2_X1 port map( A1 => n21, A2 => n25, ZN => n23);
   U34 : MUX2_X1 port map( A => n23, B => n22, S => B_isINF, Z => n24);
   U35 : NAND2_X1 port map( A1 => n26, A2 => n24, ZN => isNaN_stage1);
   U36 : NOR2_X1 port map( A1 => B_isZ, A2 => n25, ZN => n29);
   U37 : INV_X1 port map( A => n26, ZN => n27);
   U38 : NOR2_X1 port map( A1 => A_isZ, A2 => n27, ZN => n28);
   U39 : MUX2_X1 port map( A => n29, B => n28, S => B_isINF, Z => isINF_stage1)
                           ;
   U40 : XOR2_X1 port map( A => B_SIGN, B => A_SIGN, Z => SIGN_out_stage1);
   I0 : UnpackFP_0 port map( FP(31) => FP_A(31), FP(30) => FP_A(30), FP(29) => 
                           FP_A(29), FP(28) => FP_A(28), FP(27) => FP_A(27), 
                           FP(26) => FP_A(26), FP(25) => FP_A(25), FP(24) => 
                           FP_A(24), FP(23) => FP_A(23), FP(22) => FP_A(22), 
                           FP(21) => FP_A(21), FP(20) => FP_A(20), FP(19) => 
                           FP_A(19), FP(18) => FP_A(18), FP(17) => FP_A(17), 
                           FP(16) => FP_A(16), FP(15) => FP_A(15), FP(14) => 
                           FP_A(14), FP(13) => FP_A(13), FP(12) => FP_A(12), 
                           FP(11) => FP_A(11), FP(10) => FP_A(10), FP(9) => 
                           FP_A(9), FP(8) => FP_A(8), FP(7) => FP_A(7), FP(6) 
                           => FP_A(6), FP(5) => FP_A(5), FP(4) => FP_A(4), 
                           FP(3) => FP_A(3), FP(2) => FP_A(2), FP(1) => FP_A(1)
                           , FP(0) => FP_A(0), SIG(31) => n_2233, SIG(30) => 
                           n_2234, SIG(29) => n_2235, SIG(28) => n_2236, 
                           SIG(27) => n_2237, SIG(26) => n_2238, SIG(25) => 
                           n_2239, SIG(24) => n_2240, SIG(23) => A_SIG(23), 
                           SIG(22) => A_SIG(22), SIG(21) => A_SIG(21), SIG(20) 
                           => A_SIG(20), SIG(19) => A_SIG(19), SIG(18) => 
                           A_SIG(18), SIG(17) => A_SIG(17), SIG(16) => 
                           A_SIG(16), SIG(15) => A_SIG(15), SIG(14) => 
                           A_SIG(14), SIG(13) => A_SIG(13), SIG(12) => 
                           A_SIG(12), SIG(11) => A_SIG(11), SIG(10) => 
                           A_SIG(10), SIG(9) => A_SIG(9), SIG(8) => A_SIG(8), 
                           SIG(7) => A_SIG(7), SIG(6) => A_SIG(6), SIG(5) => 
                           A_SIG(5), SIG(4) => A_SIG(4), SIG(3) => A_SIG(3), 
                           SIG(2) => A_SIG(2), SIG(1) => A_SIG(1), SIG(0) => 
                           A_SIG(0), EXP(7) => A_EXP(7), EXP(6) => A_EXP(6), 
                           EXP(5) => A_EXP(5), EXP(4) => A_EXP(4), EXP(3) => 
                           A_EXP(3), EXP(2) => A_EXP(2), EXP(1) => A_EXP(1), 
                           EXP(0) => A_EXP(0), SIGN => A_SIGN, isNaN => A_isNaN
                           , isINF => A_isINF, isZ => A_isZ, isDN => n_2241);
   I1 : UnpackFP_1 port map( FP(31) => FP_B(31), FP(30) => FP_B(30), FP(29) => 
                           FP_B(29), FP(28) => FP_B(28), FP(27) => FP_B(27), 
                           FP(26) => FP_B(26), FP(25) => FP_B(25), FP(24) => 
                           FP_B(24), FP(23) => FP_B(23), FP(22) => FP_B(22), 
                           FP(21) => FP_B(21), FP(20) => FP_B(20), FP(19) => 
                           FP_B(19), FP(18) => FP_B(18), FP(17) => FP_B(17), 
                           FP(16) => FP_B(16), FP(15) => FP_B(15), FP(14) => 
                           FP_B(14), FP(13) => FP_B(13), FP(12) => FP_B(12), 
                           FP(11) => FP_B(11), FP(10) => FP_B(10), FP(9) => 
                           FP_B(9), FP(8) => FP_B(8), FP(7) => FP_B(7), FP(6) 
                           => FP_B(6), FP(5) => FP_B(5), FP(4) => FP_B(4), 
                           FP(3) => FP_B(3), FP(2) => FP_B(2), FP(1) => FP_B(1)
                           , FP(0) => FP_B(0), SIG(31) => n_2242, SIG(30) => 
                           n_2243, SIG(29) => n_2244, SIG(28) => n_2245, 
                           SIG(27) => n_2246, SIG(26) => n_2247, SIG(25) => 
                           n_2248, SIG(24) => n_2249, SIG(23) => B_SIG(23), 
                           SIG(22) => B_SIG(22), SIG(21) => B_SIG(21), SIG(20) 
                           => B_SIG(20), SIG(19) => B_SIG(19), SIG(18) => 
                           B_SIG(18), SIG(17) => B_SIG(17), SIG(16) => 
                           B_SIG(16), SIG(15) => B_SIG(15), SIG(14) => 
                           B_SIG(14), SIG(13) => B_SIG(13), SIG(12) => 
                           B_SIG(12), SIG(11) => B_SIG(11), SIG(10) => 
                           B_SIG(10), SIG(9) => B_SIG(9), SIG(8) => B_SIG(8), 
                           SIG(7) => B_SIG(7), SIG(6) => B_SIG(6), SIG(5) => 
                           B_SIG(5), SIG(4) => B_SIG(4), SIG(3) => B_SIG(3), 
                           SIG(2) => B_SIG(2), SIG(1) => B_SIG(1), SIG(0) => 
                           B_SIG(0), EXP(7) => B_EXP(7), EXP(6) => B_EXP(6), 
                           EXP(5) => B_EXP(5), EXP(4) => B_EXP(4), EXP(3) => 
                           B_EXP(3), EXP(2) => B_EXP(2), EXP(1) => B_EXP(1), 
                           EXP(0) => B_EXP(0), SIGN => B_SIGN, isNaN => B_isNaN
                           , isINF => B_isINF, isZ => B_isZ, isDN => n_2250);

end SYN_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_FPmul.all;

entity FPmul is

   port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic;  
         FP_Z : out std_logic_vector (31 downto 0));

end FPmul;

architecture SYN_pipeline of FPmul is

   component FPmul_stage4
      port( EXP_neg : in std_logic;  EXP_out_round : in std_logic_vector (7 
            downto 0);  EXP_pos, SIGN_out : in std_logic;  SIG_out_round : in 
            std_logic_vector (27 downto 0);  clk, isINF_tab, isNaN, isZ_tab : 
            in std_logic;  FP_Z : out std_logic_vector (31 downto 0));
   end component;
   
   component FPmul_stage3
      port( EXP_in : in std_logic_vector (7 downto 0);  EXP_neg_stage2, 
            EXP_pos_stage2, SIGN_out_stage2 : in std_logic;  SIG_in : in 
            std_logic_vector (27 downto 0);  clk, isINF_stage2, isNaN_stage2, 
            isZ_tab_stage2 : in std_logic;  EXP_neg : out std_logic;  
            EXP_out_round : out std_logic_vector (7 downto 0);  EXP_pos, 
            SIGN_out : out std_logic;  SIG_out_round : out std_logic_vector (27
            downto 0);  isINF_tab, isNaN, isZ_tab : out std_logic);
   end component;
   
   component FPmul_stage2
      port( A_EXP : in std_logic_vector (7 downto 0);  A_SIG : in 
            std_logic_vector (31 downto 0);  B_EXP : in std_logic_vector (7 
            downto 0);  B_SIG : in std_logic_vector (31 downto 0);  
            SIGN_out_stage1, clk, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : 
            in std_logic;  EXP_in : out std_logic_vector (7 downto 0);  
            EXP_neg_stage2, EXP_pos_stage2, SIGN_out_stage2 : out std_logic;  
            SIG_in : out std_logic_vector (27 downto 0);  isINF_stage2, 
            isNaN_stage2, isZ_tab_stage2 : out std_logic);
   end component;
   
   component FPmul_stage1
      port( FP_A, FP_B : in std_logic_vector (31 downto 0);  clk : in std_logic
            ;  A_EXP : out std_logic_vector (7 downto 0);  A_SIG : out 
            std_logic_vector (31 downto 0);  B_EXP : out std_logic_vector (7 
            downto 0);  B_SIG : out std_logic_vector (31 downto 0);  
            SIGN_out_stage1, isINF_stage1, isNaN_stage1, isZ_tab_stage1 : out 
            std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal A_EXP_7_port, A_EXP_6_port, A_EXP_5_port, A_EXP_4_port, A_EXP_3_port,
      A_EXP_2_port, A_EXP_1_port, A_EXP_0_port, A_SIG_22_port, A_SIG_21_port, 
      A_SIG_20_port, A_SIG_19_port, A_SIG_18_port, A_SIG_17_port, A_SIG_16_port
      , A_SIG_15_port, A_SIG_14_port, A_SIG_13_port, A_SIG_12_port, 
      A_SIG_11_port, A_SIG_10_port, A_SIG_9_port, A_SIG_8_port, A_SIG_7_port, 
      A_SIG_6_port, A_SIG_5_port, A_SIG_4_port, A_SIG_3_port, A_SIG_2_port, 
      A_SIG_1_port, A_SIG_0_port, B_EXP_7_port, B_EXP_6_port, B_EXP_5_port, 
      B_EXP_4_port, B_EXP_3_port, B_EXP_2_port, B_EXP_1_port, B_EXP_0_port, 
      B_SIG_22_port, B_SIG_21_port, B_SIG_20_port, B_SIG_19_port, B_SIG_18_port
      , B_SIG_17_port, B_SIG_16_port, B_SIG_15_port, B_SIG_14_port, 
      B_SIG_13_port, B_SIG_12_port, B_SIG_11_port, B_SIG_10_port, B_SIG_9_port,
      B_SIG_8_port, B_SIG_7_port, B_SIG_6_port, B_SIG_5_port, B_SIG_4_port, 
      B_SIG_3_port, B_SIG_2_port, B_SIG_1_port, B_SIG_0_port, SIGN_out_stage1, 
      isINF_stage1, isNaN_stage1, isZ_tab_stage1, EXP_in_7_port, EXP_in_6_port,
      EXP_in_5_port, EXP_in_4_port, EXP_in_3_port, EXP_in_2_port, EXP_in_1_port
      , EXP_in_0_port, EXP_neg_stage2, EXP_pos_stage2, SIGN_out_stage2, 
      SIG_in_27_port, SIG_in_26_port, SIG_in_25_port, SIG_in_24_port, 
      SIG_in_23_port, SIG_in_22_port, SIG_in_21_port, SIG_in_20_port, 
      SIG_in_19_port, SIG_in_18_port, SIG_in_17_port, SIG_in_16_port, 
      SIG_in_15_port, SIG_in_14_port, SIG_in_13_port, SIG_in_12_port, 
      SIG_in_11_port, SIG_in_10_port, SIG_in_9_port, SIG_in_8_port, 
      SIG_in_7_port, SIG_in_6_port, SIG_in_5_port, SIG_in_4_port, SIG_in_3_port
      , SIG_in_2_port, isINF_stage2, isNaN_stage2, isZ_tab_stage2, EXP_neg, 
      EXP_out_round_7_port, EXP_out_round_6_port, EXP_out_round_5_port, 
      EXP_out_round_4_port, EXP_out_round_3_port, EXP_out_round_2_port, 
      EXP_out_round_1_port, EXP_out_round_0_port, EXP_pos, SIGN_out, 
      SIG_out_round_27_port, SIG_out_round_26_port, SIG_out_round_25_port, 
      SIG_out_round_24_port, SIG_out_round_23_port, SIG_out_round_22_port, 
      SIG_out_round_21_port, SIG_out_round_20_port, SIG_out_round_19_port, 
      SIG_out_round_18_port, SIG_out_round_17_port, SIG_out_round_16_port, 
      SIG_out_round_15_port, SIG_out_round_14_port, SIG_out_round_13_port, 
      SIG_out_round_12_port, SIG_out_round_11_port, SIG_out_round_10_port, 
      SIG_out_round_9_port, SIG_out_round_8_port, SIG_out_round_7_port, 
      SIG_out_round_6_port, SIG_out_round_5_port, SIG_out_round_4_port, 
      SIG_out_round_3_port, isINF_tab, isNaN, isZ_tab, n1, n132, n88, n89, n90,
      n91, n129, n130, n131, n133, n135, n_2251, n_2252, n_2253, n_2254, n_2255
      , n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264,
      n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, 
      n_2274, n_2275 : std_logic;

begin
   
   n1 <= '0';
   n88 <= '0';
   n89 <= '0';
   n90 <= '0';
   n91 <= '0';
   MY_CLK_r_REG184_S1 : DFF_X1 port map( D => n132, CK => clk, Q => n131, QN =>
                           n_2251);
   MY_CLK_r_REG185_S2 : DFF_X1 port map( D => n131, CK => clk, Q => n130, QN =>
                           n_2252);
   MY_CLK_r_REG186_S3 : DFF_X1 port map( D => n130, CK => clk, Q => n129, QN =>
                           n_2253);
   MY_CLK_r_REG187_S4 : DFF_X1 port map( D => n129, CK => clk, Q => FP_Z(31), 
                           QN => n_2254);
   I1 : FPmul_stage1 port map( FP_A(31) => FP_A(31), FP_A(30) => FP_A(30), 
                           FP_A(29) => FP_A(29), FP_A(28) => FP_A(28), FP_A(27)
                           => FP_A(27), FP_A(26) => FP_A(26), FP_A(25) => 
                           FP_A(25), FP_A(24) => FP_A(24), FP_A(23) => FP_A(23)
                           , FP_A(22) => FP_A(22), FP_A(21) => FP_A(21), 
                           FP_A(20) => FP_A(20), FP_A(19) => FP_A(19), FP_A(18)
                           => FP_A(18), FP_A(17) => FP_A(17), FP_A(16) => 
                           FP_A(16), FP_A(15) => FP_A(15), FP_A(14) => FP_A(14)
                           , FP_A(13) => FP_A(13), FP_A(12) => FP_A(12), 
                           FP_A(11) => FP_A(11), FP_A(10) => FP_A(10), FP_A(9) 
                           => FP_A(9), FP_A(8) => FP_A(8), FP_A(7) => FP_A(7), 
                           FP_A(6) => FP_A(6), FP_A(5) => FP_A(5), FP_A(4) => 
                           FP_A(4), FP_A(3) => FP_A(3), FP_A(2) => FP_A(2), 
                           FP_A(1) => FP_A(1), FP_A(0) => FP_A(0), FP_B(31) => 
                           FP_B(31), FP_B(30) => FP_B(30), FP_B(29) => FP_B(29)
                           , FP_B(28) => FP_B(28), FP_B(27) => FP_B(27), 
                           FP_B(26) => FP_B(26), FP_B(25) => FP_B(25), FP_B(24)
                           => FP_B(24), FP_B(23) => FP_B(23), FP_B(22) => 
                           FP_B(22), FP_B(21) => FP_B(21), FP_B(20) => FP_B(20)
                           , FP_B(19) => FP_B(19), FP_B(18) => FP_B(18), 
                           FP_B(17) => FP_B(17), FP_B(16) => FP_B(16), FP_B(15)
                           => FP_B(15), FP_B(14) => FP_B(14), FP_B(13) => 
                           FP_B(13), FP_B(12) => FP_B(12), FP_B(11) => FP_B(11)
                           , FP_B(10) => FP_B(10), FP_B(9) => FP_B(9), FP_B(8) 
                           => FP_B(8), FP_B(7) => FP_B(7), FP_B(6) => FP_B(6), 
                           FP_B(5) => FP_B(5), FP_B(4) => FP_B(4), FP_B(3) => 
                           FP_B(3), FP_B(2) => FP_B(2), FP_B(1) => FP_B(1), 
                           FP_B(0) => FP_B(0), clk => clk, A_EXP(7) => 
                           A_EXP_7_port, A_EXP(6) => A_EXP_6_port, A_EXP(5) => 
                           A_EXP_5_port, A_EXP(4) => A_EXP_4_port, A_EXP(3) => 
                           A_EXP_3_port, A_EXP(2) => A_EXP_2_port, A_EXP(1) => 
                           A_EXP_1_port, A_EXP(0) => A_EXP_0_port, A_SIG(31) =>
                           n_2255, A_SIG(30) => n_2256, A_SIG(29) => n_2257, 
                           A_SIG(28) => n_2258, A_SIG(27) => n_2259, A_SIG(26) 
                           => n_2260, A_SIG(25) => n_2261, A_SIG(24) => n_2262,
                           A_SIG(23) => n135, A_SIG(22) => A_SIG_22_port, 
                           A_SIG(21) => A_SIG_21_port, A_SIG(20) => 
                           A_SIG_20_port, A_SIG(19) => A_SIG_19_port, A_SIG(18)
                           => A_SIG_18_port, A_SIG(17) => A_SIG_17_port, 
                           A_SIG(16) => A_SIG_16_port, A_SIG(15) => 
                           A_SIG_15_port, A_SIG(14) => A_SIG_14_port, A_SIG(13)
                           => A_SIG_13_port, A_SIG(12) => A_SIG_12_port, 
                           A_SIG(11) => A_SIG_11_port, A_SIG(10) => 
                           A_SIG_10_port, A_SIG(9) => A_SIG_9_port, A_SIG(8) =>
                           A_SIG_8_port, A_SIG(7) => A_SIG_7_port, A_SIG(6) => 
                           A_SIG_6_port, A_SIG(5) => A_SIG_5_port, A_SIG(4) => 
                           A_SIG_4_port, A_SIG(3) => A_SIG_3_port, A_SIG(2) => 
                           A_SIG_2_port, A_SIG(1) => A_SIG_1_port, A_SIG(0) => 
                           A_SIG_0_port, B_EXP(7) => B_EXP_7_port, B_EXP(6) => 
                           B_EXP_6_port, B_EXP(5) => B_EXP_5_port, B_EXP(4) => 
                           B_EXP_4_port, B_EXP(3) => B_EXP_3_port, B_EXP(2) => 
                           B_EXP_2_port, B_EXP(1) => B_EXP_1_port, B_EXP(0) => 
                           B_EXP_0_port, B_SIG(31) => n_2263, B_SIG(30) => 
                           n_2264, B_SIG(29) => n_2265, B_SIG(28) => n_2266, 
                           B_SIG(27) => n_2267, B_SIG(26) => n_2268, B_SIG(25) 
                           => n_2269, B_SIG(24) => n_2270, B_SIG(23) => n133, 
                           B_SIG(22) => B_SIG_22_port, B_SIG(21) => 
                           B_SIG_21_port, B_SIG(20) => B_SIG_20_port, B_SIG(19)
                           => B_SIG_19_port, B_SIG(18) => B_SIG_18_port, 
                           B_SIG(17) => B_SIG_17_port, B_SIG(16) => 
                           B_SIG_16_port, B_SIG(15) => B_SIG_15_port, B_SIG(14)
                           => B_SIG_14_port, B_SIG(13) => B_SIG_13_port, 
                           B_SIG(12) => B_SIG_12_port, B_SIG(11) => 
                           B_SIG_11_port, B_SIG(10) => B_SIG_10_port, B_SIG(9) 
                           => B_SIG_9_port, B_SIG(8) => B_SIG_8_port, B_SIG(7) 
                           => B_SIG_7_port, B_SIG(6) => B_SIG_6_port, B_SIG(5) 
                           => B_SIG_5_port, B_SIG(4) => B_SIG_4_port, B_SIG(3) 
                           => B_SIG_3_port, B_SIG(2) => B_SIG_2_port, B_SIG(1) 
                           => B_SIG_1_port, B_SIG(0) => B_SIG_0_port, 
                           SIGN_out_stage1 => SIGN_out_stage1, isINF_stage1 => 
                           isINF_stage1, isNaN_stage1 => isNaN_stage1, 
                           isZ_tab_stage1 => isZ_tab_stage1);
   I2 : FPmul_stage2 port map( A_EXP(7) => A_EXP_7_port, A_EXP(6) => 
                           A_EXP_6_port, A_EXP(5) => A_EXP_5_port, A_EXP(4) => 
                           A_EXP_4_port, A_EXP(3) => A_EXP_3_port, A_EXP(2) => 
                           A_EXP_2_port, A_EXP(1) => A_EXP_1_port, A_EXP(0) => 
                           A_EXP_0_port, A_SIG(31) => n1, A_SIG(30) => n1, 
                           A_SIG(29) => n1, A_SIG(28) => n1, A_SIG(27) => n1, 
                           A_SIG(26) => n1, A_SIG(25) => n1, A_SIG(24) => n1, 
                           A_SIG(23) => n135, A_SIG(22) => A_SIG_22_port, 
                           A_SIG(21) => A_SIG_21_port, A_SIG(20) => 
                           A_SIG_20_port, A_SIG(19) => A_SIG_19_port, A_SIG(18)
                           => A_SIG_18_port, A_SIG(17) => A_SIG_17_port, 
                           A_SIG(16) => A_SIG_16_port, A_SIG(15) => 
                           A_SIG_15_port, A_SIG(14) => A_SIG_14_port, A_SIG(13)
                           => A_SIG_13_port, A_SIG(12) => A_SIG_12_port, 
                           A_SIG(11) => A_SIG_11_port, A_SIG(10) => 
                           A_SIG_10_port, A_SIG(9) => A_SIG_9_port, A_SIG(8) =>
                           A_SIG_8_port, A_SIG(7) => A_SIG_7_port, A_SIG(6) => 
                           A_SIG_6_port, A_SIG(5) => A_SIG_5_port, A_SIG(4) => 
                           A_SIG_4_port, A_SIG(3) => A_SIG_3_port, A_SIG(2) => 
                           A_SIG_2_port, A_SIG(1) => A_SIG_1_port, A_SIG(0) => 
                           A_SIG_0_port, B_EXP(7) => B_EXP_7_port, B_EXP(6) => 
                           B_EXP_6_port, B_EXP(5) => B_EXP_5_port, B_EXP(4) => 
                           B_EXP_4_port, B_EXP(3) => B_EXP_3_port, B_EXP(2) => 
                           B_EXP_2_port, B_EXP(1) => B_EXP_1_port, B_EXP(0) => 
                           B_EXP_0_port, B_SIG(31) => n1, B_SIG(30) => n1, 
                           B_SIG(29) => n1, B_SIG(28) => n1, B_SIG(27) => n1, 
                           B_SIG(26) => n1, B_SIG(25) => n1, B_SIG(24) => n1, 
                           B_SIG(23) => n133, B_SIG(22) => B_SIG_22_port, 
                           B_SIG(21) => B_SIG_21_port, B_SIG(20) => 
                           B_SIG_20_port, B_SIG(19) => B_SIG_19_port, B_SIG(18)
                           => B_SIG_18_port, B_SIG(17) => B_SIG_17_port, 
                           B_SIG(16) => B_SIG_16_port, B_SIG(15) => 
                           B_SIG_15_port, B_SIG(14) => B_SIG_14_port, B_SIG(13)
                           => B_SIG_13_port, B_SIG(12) => B_SIG_12_port, 
                           B_SIG(11) => B_SIG_11_port, B_SIG(10) => 
                           B_SIG_10_port, B_SIG(9) => B_SIG_9_port, B_SIG(8) =>
                           B_SIG_8_port, B_SIG(7) => B_SIG_7_port, B_SIG(6) => 
                           B_SIG_6_port, B_SIG(5) => B_SIG_5_port, B_SIG(4) => 
                           B_SIG_4_port, B_SIG(3) => B_SIG_3_port, B_SIG(2) => 
                           B_SIG_2_port, B_SIG(1) => B_SIG_1_port, B_SIG(0) => 
                           B_SIG_0_port, SIGN_out_stage1 => SIGN_out_stage1, 
                           clk => clk, isINF_stage1 => isINF_stage1, 
                           isNaN_stage1 => isNaN_stage1, isZ_tab_stage1 => 
                           isZ_tab_stage1, EXP_in(7) => EXP_in_7_port, 
                           EXP_in(6) => EXP_in_6_port, EXP_in(5) => 
                           EXP_in_5_port, EXP_in(4) => EXP_in_4_port, EXP_in(3)
                           => EXP_in_3_port, EXP_in(2) => EXP_in_2_port, 
                           EXP_in(1) => EXP_in_1_port, EXP_in(0) => 
                           EXP_in_0_port, EXP_neg_stage2 => EXP_neg_stage2, 
                           EXP_pos_stage2 => EXP_pos_stage2, SIGN_out_stage2 =>
                           SIGN_out_stage2, SIG_in(27) => SIG_in_27_port, 
                           SIG_in(26) => SIG_in_26_port, SIG_in(25) => 
                           SIG_in_25_port, SIG_in(24) => SIG_in_24_port, 
                           SIG_in(23) => SIG_in_23_port, SIG_in(22) => 
                           SIG_in_22_port, SIG_in(21) => SIG_in_21_port, 
                           SIG_in(20) => SIG_in_20_port, SIG_in(19) => 
                           SIG_in_19_port, SIG_in(18) => SIG_in_18_port, 
                           SIG_in(17) => SIG_in_17_port, SIG_in(16) => 
                           SIG_in_16_port, SIG_in(15) => SIG_in_15_port, 
                           SIG_in(14) => SIG_in_14_port, SIG_in(13) => 
                           SIG_in_13_port, SIG_in(12) => SIG_in_12_port, 
                           SIG_in(11) => SIG_in_11_port, SIG_in(10) => 
                           SIG_in_10_port, SIG_in(9) => SIG_in_9_port, 
                           SIG_in(8) => SIG_in_8_port, SIG_in(7) => 
                           SIG_in_7_port, SIG_in(6) => SIG_in_6_port, SIG_in(5)
                           => SIG_in_5_port, SIG_in(4) => SIG_in_4_port, 
                           SIG_in(3) => SIG_in_3_port, SIG_in(2) => 
                           SIG_in_2_port, SIG_in(1) => n_2271, SIG_in(0) => 
                           n_2272, isINF_stage2 => isINF_stage2, isNaN_stage2 
                           => isNaN_stage2, isZ_tab_stage2 => isZ_tab_stage2);
   I3 : FPmul_stage3 port map( EXP_in(7) => EXP_in_7_port, EXP_in(6) => 
                           EXP_in_6_port, EXP_in(5) => EXP_in_5_port, EXP_in(4)
                           => EXP_in_4_port, EXP_in(3) => EXP_in_3_port, 
                           EXP_in(2) => EXP_in_2_port, EXP_in(1) => 
                           EXP_in_1_port, EXP_in(0) => EXP_in_0_port, 
                           EXP_neg_stage2 => EXP_neg_stage2, EXP_pos_stage2 => 
                           EXP_pos_stage2, SIGN_out_stage2 => SIGN_out_stage2, 
                           SIG_in(27) => SIG_in_27_port, SIG_in(26) => 
                           SIG_in_26_port, SIG_in(25) => SIG_in_25_port, 
                           SIG_in(24) => SIG_in_24_port, SIG_in(23) => 
                           SIG_in_23_port, SIG_in(22) => SIG_in_22_port, 
                           SIG_in(21) => SIG_in_21_port, SIG_in(20) => 
                           SIG_in_20_port, SIG_in(19) => SIG_in_19_port, 
                           SIG_in(18) => SIG_in_18_port, SIG_in(17) => 
                           SIG_in_17_port, SIG_in(16) => SIG_in_16_port, 
                           SIG_in(15) => SIG_in_15_port, SIG_in(14) => 
                           SIG_in_14_port, SIG_in(13) => SIG_in_13_port, 
                           SIG_in(12) => SIG_in_12_port, SIG_in(11) => 
                           SIG_in_11_port, SIG_in(10) => SIG_in_10_port, 
                           SIG_in(9) => SIG_in_9_port, SIG_in(8) => 
                           SIG_in_8_port, SIG_in(7) => SIG_in_7_port, SIG_in(6)
                           => SIG_in_6_port, SIG_in(5) => SIG_in_5_port, 
                           SIG_in(4) => SIG_in_4_port, SIG_in(3) => 
                           SIG_in_3_port, SIG_in(2) => SIG_in_2_port, SIG_in(1)
                           => n88, SIG_in(0) => n89, clk => clk, isINF_stage2 
                           => isINF_stage2, isNaN_stage2 => isNaN_stage2, 
                           isZ_tab_stage2 => isZ_tab_stage2, EXP_neg => EXP_neg
                           , EXP_out_round(7) => EXP_out_round_7_port, 
                           EXP_out_round(6) => EXP_out_round_6_port, 
                           EXP_out_round(5) => EXP_out_round_5_port, 
                           EXP_out_round(4) => EXP_out_round_4_port, 
                           EXP_out_round(3) => EXP_out_round_3_port, 
                           EXP_out_round(2) => EXP_out_round_2_port, 
                           EXP_out_round(1) => EXP_out_round_1_port, 
                           EXP_out_round(0) => EXP_out_round_0_port, EXP_pos =>
                           EXP_pos, SIGN_out => SIGN_out, SIG_out_round(27) => 
                           SIG_out_round_27_port, SIG_out_round(26) => 
                           SIG_out_round_26_port, SIG_out_round(25) => 
                           SIG_out_round_25_port, SIG_out_round(24) => 
                           SIG_out_round_24_port, SIG_out_round(23) => 
                           SIG_out_round_23_port, SIG_out_round(22) => 
                           SIG_out_round_22_port, SIG_out_round(21) => 
                           SIG_out_round_21_port, SIG_out_round(20) => 
                           SIG_out_round_20_port, SIG_out_round(19) => 
                           SIG_out_round_19_port, SIG_out_round(18) => 
                           SIG_out_round_18_port, SIG_out_round(17) => 
                           SIG_out_round_17_port, SIG_out_round(16) => 
                           SIG_out_round_16_port, SIG_out_round(15) => 
                           SIG_out_round_15_port, SIG_out_round(14) => 
                           SIG_out_round_14_port, SIG_out_round(13) => 
                           SIG_out_round_13_port, SIG_out_round(12) => 
                           SIG_out_round_12_port, SIG_out_round(11) => 
                           SIG_out_round_11_port, SIG_out_round(10) => 
                           SIG_out_round_10_port, SIG_out_round(9) => 
                           SIG_out_round_9_port, SIG_out_round(8) => 
                           SIG_out_round_8_port, SIG_out_round(7) => 
                           SIG_out_round_7_port, SIG_out_round(6) => 
                           SIG_out_round_6_port, SIG_out_round(5) => 
                           SIG_out_round_5_port, SIG_out_round(4) => 
                           SIG_out_round_4_port, SIG_out_round(3) => 
                           SIG_out_round_3_port, SIG_out_round(2) => n_2273, 
                           SIG_out_round(1) => n_2274, SIG_out_round(0) => 
                           n_2275, isINF_tab => isINF_tab, isNaN => isNaN, 
                           isZ_tab => isZ_tab);
   I4 : FPmul_stage4 port map( EXP_neg => EXP_neg, EXP_out_round(7) => 
                           EXP_out_round_7_port, EXP_out_round(6) => 
                           EXP_out_round_6_port, EXP_out_round(5) => 
                           EXP_out_round_5_port, EXP_out_round(4) => 
                           EXP_out_round_4_port, EXP_out_round(3) => 
                           EXP_out_round_3_port, EXP_out_round(2) => 
                           EXP_out_round_2_port, EXP_out_round(1) => 
                           EXP_out_round_1_port, EXP_out_round(0) => 
                           EXP_out_round_0_port, EXP_pos => EXP_pos, SIGN_out 
                           => SIGN_out, SIG_out_round(27) => 
                           SIG_out_round_27_port, SIG_out_round(26) => 
                           SIG_out_round_26_port, SIG_out_round(25) => 
                           SIG_out_round_25_port, SIG_out_round(24) => 
                           SIG_out_round_24_port, SIG_out_round(23) => 
                           SIG_out_round_23_port, SIG_out_round(22) => 
                           SIG_out_round_22_port, SIG_out_round(21) => 
                           SIG_out_round_21_port, SIG_out_round(20) => 
                           SIG_out_round_20_port, SIG_out_round(19) => 
                           SIG_out_round_19_port, SIG_out_round(18) => 
                           SIG_out_round_18_port, SIG_out_round(17) => 
                           SIG_out_round_17_port, SIG_out_round(16) => 
                           SIG_out_round_16_port, SIG_out_round(15) => 
                           SIG_out_round_15_port, SIG_out_round(14) => 
                           SIG_out_round_14_port, SIG_out_round(13) => 
                           SIG_out_round_13_port, SIG_out_round(12) => 
                           SIG_out_round_12_port, SIG_out_round(11) => 
                           SIG_out_round_11_port, SIG_out_round(10) => 
                           SIG_out_round_10_port, SIG_out_round(9) => 
                           SIG_out_round_9_port, SIG_out_round(8) => 
                           SIG_out_round_8_port, SIG_out_round(7) => 
                           SIG_out_round_7_port, SIG_out_round(6) => 
                           SIG_out_round_6_port, SIG_out_round(5) => 
                           SIG_out_round_5_port, SIG_out_round(4) => 
                           SIG_out_round_4_port, SIG_out_round(3) => 
                           SIG_out_round_3_port, SIG_out_round(2) => n1, 
                           SIG_out_round(1) => n90, SIG_out_round(0) => n91, 
                           clk => clk, isINF_tab => isINF_tab, isNaN => isNaN, 
                           isZ_tab => isZ_tab, FP_Z(31) => n132, FP_Z(30) => 
                           FP_Z(30), FP_Z(29) => FP_Z(29), FP_Z(28) => FP_Z(28)
                           , FP_Z(27) => FP_Z(27), FP_Z(26) => FP_Z(26), 
                           FP_Z(25) => FP_Z(25), FP_Z(24) => FP_Z(24), FP_Z(23)
                           => FP_Z(23), FP_Z(22) => FP_Z(22), FP_Z(21) => 
                           FP_Z(21), FP_Z(20) => FP_Z(20), FP_Z(19) => FP_Z(19)
                           , FP_Z(18) => FP_Z(18), FP_Z(17) => FP_Z(17), 
                           FP_Z(16) => FP_Z(16), FP_Z(15) => FP_Z(15), FP_Z(14)
                           => FP_Z(14), FP_Z(13) => FP_Z(13), FP_Z(12) => 
                           FP_Z(12), FP_Z(11) => FP_Z(11), FP_Z(10) => FP_Z(10)
                           , FP_Z(9) => FP_Z(9), FP_Z(8) => FP_Z(8), FP_Z(7) =>
                           FP_Z(7), FP_Z(6) => FP_Z(6), FP_Z(5) => FP_Z(5), 
                           FP_Z(4) => FP_Z(4), FP_Z(3) => FP_Z(3), FP_Z(2) => 
                           FP_Z(2), FP_Z(1) => FP_Z(1), FP_Z(0) => FP_Z(0));

end SYN_pipeline;
