package pkgfla is
	constant nb : integer := 14;
	constant r : integer := 5;
	constant nb_w : integer := 17;
	constant nb_a : integer := 22;
end pkgfla;
