package my_pkg is

	constant n_levels : integer := 7;

  type rows_type is array (7 downto 0) of integer;
  constant row, col_start, col_end, num_start, num_end : rows_type;
  
end my_pkg;

package body my_pkg is 

  constant row        : rows_type := (17,13, 9, 6, 4, 3, 2, 2);
  constant col_start  : rows_type := (24,16,10, 6, 4, 2, 0, 0);
  constant col_end    : rows_type := (42,50,56,60,62,64, 0, 0);

  constant num_start  : rows_type := ( 0, 8,16,22,26,28, 0, 0);
  constant num_end    : rows_type := ( 8, 8, 6, 4, 2, 2, 0, 0);

end my_pkg;
